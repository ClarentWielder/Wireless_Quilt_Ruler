PK   F�X�pǿ�  �C     cirkitFile.json�Qo�6��ʠ��I���u�C�(�=āA[t#̑<YN����Q�dǒM��a�F�ݑ�;�Y�kT�gSΗUm�Ϧ�U�P1�u����V2�6E9o���Zo��W��6�7f���6Ui�fNY��b�\dl�US�36%�d���Z�9�n�&�V�8u�SOp��.p�)N=��Cʋt��ҜL��U��JM�r%�iB�XR��F۱#K��fd��;�v�ĝ"y�H�)�x�D�fH}��G���s�s�-G��Rw:/�q��Rw9/�q��Rw8/�q���{�y� F;�<���c���� �V��	f�'��>��.�l~���~ti�ZW52��~&���� VX+I+<��J�JĊ+�Ҋ
C] x��K��K��K� L�L� L�0Le3a(f�u)#Øi)6|���$��|s� V�:�of��Uw��SX��L����H�F�N]s��.�a�~xg|��>��6�1�į4���kd⇷XI�X�A�� V� V� Vd+*u��C/�/�/0C0�0�01C1C1�J�w⇷f.W�;��[��Nމ��Ug�N��V���w���@�����y�����į4ߚ���y��n�$z)j��o�V>�ۼ��sSG7������a�yҊ�p0#K\���p���Á��<U�]�C<��I�gP<��	 ��O �~hR�]绢���Z�����9���#+J�>C�'H}��H���9��|��]6�1�}p���'�O��b	�XD)�Q���Ճ(k K����8F�-���|�z�Q�+A��7��0��Ļ����qػ�����_@ؔ�/�׃(x��^������^��!?�����Dx��ȁ����폰?�TCf�-d��	�$Q
��)HS� OA����U �5�&/���;P�n��}��j�K�����cQ��*�sE�و,�����'��Yj�[��^���3��?L��x�����w�};�J�]	8�^����|Q�B���j�.�M��xO���o��zuMwu�1uS�6%�7Ȏ�m��j�S�'���I���;�b��2veaG��o����S��5ݬ�zkl���_�m�X���6���r��wƮ�I���^6��ԗF?��K�W��h~�-��ؕ�g�L�mѸ���B�*#L$\�O:a���W�o���o��(Y,�$�f��H)nI��t�u�0�9Y�aݞ|�� e�@��r��
ד���.my�lD��.�������j�b�2;�{!��M�8s2�DX+"I�BAF�$ݯw��U�ک�F9q&"{��-;|�T���Tꤘ��)�Ÿ�I>��OI���'T�������X;)*�a������ڇ���^֎KG����<LolX�n����Hw���H`?�۽�q9[αX��p�Cr�����W�|nvyQu��8�����ȕ$.%�?D.
�K�R�&��}���h���T�DMW#�)Y�)�DjnRj��+Xy�s��2�Rb)���)��䡣u*�2խ��pnd��!��C��+�uƝ����A͵�D���3"zI����N���3�S��7b�f1͒��T6"g�T�x�B��1aRp�/���F�T��7ӊ%	S�h2N2�0z4�1�뒥�wM�bv/u�9!�ve�6�c��sۍ^�Н�XH�B�K�7��Is*��M����`���}?��^>��C� �զi�)�˟���Y��͢���-�Y4�Y��usW����zw22�hʯ�p�j��9�Ԭ����nSes��Gg�u6�E�o~Z�A�g��zs���8����9.L�2(��q��T��D�s�����E���X�����'�O�.|�T�">�R#`�����[)F!��E/����E8İ���Mڐ(2�E����B�(��K^��<�b��|+�_�E)?�>��Й�0@�K�A"� R�"AR����.�F��)�:��O�f����)?�>g=�z�T#���z�i�Q7�.lUcS;���]����-���C�tۘ����1c��_PK   F�X����V5 GH /   images/553717b1-fb1f-43bb-91a8-4009c3c39665.pngl{P\A����A��;�wwww�����������[�����(�^1L���=����f�~H"���  $i)1%  j  σ�����.��"�*��X�0��pR��  q����RE4��"��lo��n�d
pwwg���v66t0e�w2O��� � �ž�xd���{(�/<�5u�|u'صb�ĕc����FG��B���r�g�+q�u�11U���-l88�U�cS��z��2�+W�#
X������x�������7�<����;[��TR�n.?	�+��H ��Ve�|jL����}9̃�B�B���0��{�v���k�ч"�  k������s!���4X�2��:�����!�I���"���%�fe������2��w�����
������Љ4x� ��Rw��[��W���>�el����$�>�	Lǭ��E��p(�q��N����gm�A0`�;ʰ�G�
m%kC�20��_���c�k�D�;�\ǦCx�
���@�M���]�\ ���&#��:�ی�U�]� �L��~�Q��s���2����@��p��Ou���	�G84��8��w�
�E8�)��k�!`�n��x�$�=���P]4�5J�)%�Ԁ'�c�j�/��<������z�Ĥ13��i3��4���I� lq ��VE�5g�Y�_4^}�g���s�n;TQ��B`W�ֿɜ81G$-�C������n~�����z!Z̴��Rwl*���E�C�Q����ț>�q�!N�C�'AYx�o�+D�V�w��B�k�rq	zy!_��V ���0O?T��-��ҳ���9uj�d�
�х��Q���+�������T�lj��Q�"-��4U(�˜:.Qk$w���%��Bc����>�r���ηʟ,B�	�ؓ�����ey?�Tn'I�$��qj��S�Ggg����#-5`op]� �	��edwzϕ��ęUHhh2NNl444X8�o�>��9j���c8�؟����vv��l�����55����!cbB���<:�GF���M�Ρ���#Dbʎ��wB#"B�����p����iimUTW}{�I��P��R�����vHv&2���ۉ?�3,V, �*��p��Q$�����������s�o�b�$J:�V�Q���8�)}�������Z�$}������/�IH��
�`��-/CxS-((/�:x����qG��
�z�j��f�
+�7�:|��OAs*O*�\�Z�{��p����B! ��$\�Ł !,�ߐZX� �XֆOI�܍��*��fJ%���g��<�t�����!&�ha�ۛ��iPâ�Kna�x?G��BH�̊~�Z�7A���I{�F�>Ng"���v8���͸�&�A��in/�Ǧ�����r��?���$#�����.8�����̴�g�5Fӑ�ۭ�D�Z�6�I��\�An�� �Y�+>�ڗ������R2̎mj�� ���)0�gʛ��111�Z�6��������;��ls@�fJ���l����Si�A�<Ԅ���Ǫ�`�{��k�~��b�x�����m��V�sf� ����F��xzF~��]^*� ��O����:�25�Kg�����5��QK��#��zp" La�뛖���ҷ�k��D@JQc��e��=Q?yЅ��w�� 8����V�H�j���: R{x#�ҁ��V]i���ߐ
P�Z��)^ݸ��x��0ftj�%��(���	#� �-�]�!>��0�4i$�*�Ξ}�3I�%�@R��%�#)@5�#�z.P�J8[%a$�9G�
�NO?xwfhZ���ŪN�l�"�s��8�e9�'�������Z4v��VX-Ѽ�ݷhGU��a�W�$���]��L5��q���p�T�|x�^pq+��f�n^mpֳ��@�3�Ǧ�����X���RW�a�(q8��T	}G�v���27��s6�� �;��v�V��?���>ާN�ԆX���f��� ?vP�ӧ�+K�Q:5W�lB*j��N���F�\�c
�Wh;�"����۟�Դ�\�]�XJ�8 Q	�/ej�����Qj2�4����������]jA�	:5uE���R��e"V��ujRK��c<���ql'Y�F��'Rͧc��5���h�a���u�H}p��*�?!��ZrB4{,9o��>��8���c�V��}����KԶ:��S��Ծ>y��T� ��˺�.������)]��p��{ �������n���)�Ҥ�Äez�b3)�y�/6����y�t.��_Hg�����4p)�8`���Z��������IS�������⇢��y��^&���y��?4�.D ��	}Y,�e���i����̕��Qfff.՚�4خ��}}Xw��.��1rG D�	�VԨv��WB���?H��,�+(��K	�-��`$*�U�cL�U�jP�#�x���������\����0=0�/�;�<�;���ŞUL�n��ji�h�I*K��l�Pe-6g�a��Yx�E�pO�4;�
��v8l���G-��xȁ�1P͇��<�w*��#̋Ϭ�1�(�l�l��~�B9SugpKԳ��I	y�>d��'ׯ�y�e��H�=p��[�;�e��d\K����
��!��.���
l\�
�V�� �r����;��^J���g��%��] V��bcbc��
]<|#�����ڤMf�X�[|Xx�;n������o=���-Jӛ<$'ˮ�s�}�9�m�P�ʎ.��=�A�ro\.o+I%����B�j��\���I	���Qv_2�Skkٔ�?�)T�dЋA�g�KВ7eq�䢍_��R��R���������>�'\��}镥��w��h|��Wv��P�{� �^�Db����@ίyZ[_��HH�Ɨ��. R�	YS�*�#H�K���tSԭJ���lN{�37���ҫ���F���rv�*��o�/������Uƃ�6+u�W�i
zz����osKUn?uiHl�5���=��"`�wu���A�(��
|'�
����Ӟ��#c���c�F;��͘�l?����(̐���������t��@@k+��X��Ϭbaa����}�ڰ"�B�*M<��F1�qI���!8Ƞ��_��9��&��k����&�Ɨ�rj��(���I��No�s����dO��S��nJ8�� p���>��ʂ�҈≟�&�W���6��}s���&]N: q7�k�?_� ��Kq=R��5��+�����s�� t���K����j��5l8�X�	{^���-,��-�_`��"z)� |;4y�lhh/'%.�Pm_�ϊ�7
�^Pqty���k���Vw�W|>�&��G�%��=Q�e�x`�cC���ѩ�\����W
��s�3y��GaDZ(���"���Q4� �<C���<e�=�X�&�GNoBeOz_��
x?�mhp��~xx ��gf�����w�O�	N���?�oU6���&g`@bMEd``@�짦��%�LA��0K �����Ӷ
@¡x�m�Q�/$��yu4Tf�A;ww�������ȝ��II9ee����~�2�d�RՀ ������e 	c<W�-��7��ЬS�Q>��4���}}(��|2���R��?�G�(��;x|8*ql�q{xU�I��e��o�P)f�g`"�He�����5�9���sQBd�̓�i�D�`�KĚ*�v�E�����v_B��v'�_��Uپ�$/X�,)�7�4k	TQ�]\(��ۆ�M3��v��h���}^O�z��u.��bY���Wu0��c��BZ�{��|B��\Us�G��I�ن�m>y�JF�}��wu��>���m��yx��[
Z�L~x I�>{�?#�� -
������x't� ���e�3?1�v<�|�Ї�J�����(EM���ȈS��o
� 6�wo�V��g�@���k���;�����N$���id�^f���w}�%�2ڬ�-��c���ԭ�.�60y���xW�����ƈd�8��ۣ{/Я��U��U=�l����r-���M�@��ю�F�6�V0�d�V��A�gք��+a�k�͚6���x}��d;� wS]2X=���s�w�tՀ��"UӪui�H��AL�{	LS��[Ǜ�p�	����H�'q�.��SR�н�۹0]v\����t��b�������ړQ�j�z˩��K���;^�gP_�t�����n��&cv'8M�?�6����"�Lȭ�����)�L�_mU1j1oͼ���ē��l|�4�9�	�2�K�<[�M�̖0`0cb�֕��m�w�~��'� ���KN>��h`S{Z�N�`�e�]d�	xtW����j�y����\��2�>�#�ı"n�?� H ���p�ȏ� �.ä�OXEzC5��>n��%�y�_����}�=�3hL:80;[�G QAp��ӓ�B��F��E�m�؅6sdV6���P���޸Ə�tҚ"/[�Tʺ=�~� g���'�C����)}��`knq{VF�r["�Gp"�Т,)G�ό�ZX�I�o����%~li�h�s�ki�=YnN��M��ˊJ �g��݌"�[�D� ̙�O7��<��(�gJ���o��0����,y�UnI֖I���Z��>�˅w� ��/K�EG�KK��>�E����F���M6�c��N&��_ ��UMa�	��'d�����y����(�!ۊ8�_6M�!�]���,R�kM:|�Y�(1�ʵB��)��d�v�rDA��<�}vH���>1�`���g�	��rh{XeN��huc`Ǐb�G����-�_����E�
w��WJ�	��������4�dkee��vR��t���i/l�|��������f�����B������q,�m��o����ɠ?�i��/�v�����3G��
����CP[��x�%%��u���,.�O�?5�QKT������wզn5�ܖ��XY�>�EZ�/,��̢j[����C�rҧ�ʕ��4�!j�"�j�A}���uK�:�v�Y�t5��}�ZY ��Hidr�9h^�IS�Xj��R�3�x��h���Ƭ�%��=��C+Sx~rq\o�.��ͪޣ��:���|��3;m�XnR�}�V���������8���Q��1#�R�|�J���n^J�����y�"	�ţ�DD��Ibw���oF$t��@�ւ���E��`RW�%%zs���fT,�evDD�Dr	���q�k�r��v�D���:�:�
�˭ǃ��T��
G��!�to����Õ����i�����,�]z'�%�
5��_�
ixOO���K�Y+Z�A����<E"��h`h򸰩�l��B�1�vd|vvl\\��f��]��5�Z�Nx.Y����>��պ�it�r������|�������Ia���XO>�/'tC&� �w||,���t���z���� �"���zW�;�PPj�q������������ؠw@����W����{�o�8�d؟{V��9
 ��Ь,=���@ ̺ ���[^�f�ʋ�W]NG��ye{;�v�]�B�6:z`4���@t����T��"�v�Mw��ڭ�Hڻ��n��z��Gp��D\�+�*�7/o����H�BI���)Y�r�ƈ*Z��S��}fl����� ~zF�lDo����ȋ�߫&E{��^���Op�&]�o�v�J���ﱮ�k�_��V��[���H�|�,R	uR����������$����#�D��y��޵L�\�������F�E��I�Z�F����M��C�k�d�c��F�tXn��J�I�:��"��,�kHRA~_q���`q�D0TT���lD/X���J[9W���	�*��P6���7u��Ԋ��~�5�o���I�sb���n|%�G��G��^9C�\�P��4[h?�PQ�,!ٳ�t���)U�`���EM]RRRa�!�:��"�ٽ!��<A�t[ �T�T�����ʹ��wo�
��N�6L�r6�D�p1����v	�?s*�s���r��;�_ˑ�t��e�Q�@Z�YYטd�t��\u3V|�S����N����lP���0K��Ҧ�a�	N�.#6vp��*@�Z�"QM�F�"+�����E�� ���^���(b_	�ϑ��1޺r��B4r\4��l�n*r��'x���':g%��r���c!brwD��#�E��f��l�_���Mp����]�u�s��P=�VN�ܧ���SO� �^0;�G��N@��h0 �PD33_�afh9x��)p�/�ZhX$ \Y�Ǌ5�>�����t�[�}�Γ�+*��s��?]$M�KH����F���Ka�D��hb@��W �h��R�PR��]}5���������	yZo��Egq�&�b�tPC~�Kmuz^�b>ݾ#|8����	ž㹐A�C�r
Qf� ��x��AH�������}(���x���q��L��sG�{��� 2h����l٘�E��9}��j����"����:׿Mu��!�{��8�� a�քV����B{zoʁ��P�{��:�Fɗя@ex(]��:FG��,�m��L�s3Q����NkmaQ���WA����'Sy���y����D63)�i�T�1n�r���T�+�)
q�C�]�嬑��KIgX:�[�m�1q�{;��o�*%���u��O����q�����?�s��̧�ǎʅ}�=�x\�>��?:G=M=�mz���N�h Zq�Z���H�٩�Yq}�5Šb��#�����OD�$%�.s�}�ι|lQ�5f�D�l�%j�d��� �`���ǁ;��pf�ĸ]4��3����K�h�_��i���SĆ���lyrU��9Z�������$L�����	p7�$B�Dl>n�~w�MӜ5��P�fM�K�vj/-��
J=��m��0!A!9^ ���'C�٪��&Ey�l΄j��v�, X\N���R���q��U���D�X��l��w=�q��ƺfHF;Ǐ�G��=�͛>[Kh)-|$���xd�߀�`�oh�6��q51�h�`�$��!��jNF��_�}7��D��CIo��`k�~�_�֜"�
�}d:���Y�ZфN���ļ�գ�e�/4���)iOM�C�okH|Ǉ	!�
�r�#�^����(����z�Y�.P?�Iď�[���j+�:��$��G����9��屙c�%�=ah�
���׿�`H|P�~�,�!�ۣ�?���y~�#ԃ�l�Eg��"�NG��'#W��]�1����t�qsڔ�w4�2m��ȣ�����4d�e����;��9\k�'�f�	�E1��_�P� M�8�w�� ���.t� 10\(^�oKzQZÄL��T��\�ȴq�~o>���aaaU+K����oO�tIJr�b6r�=��x��@���i�?��_�Wy:�Syě���)��U�N[TY�R��MKz����n`�C}�۔(��/�K����?o5I�B��������%sV����c�N{k���vP�O���n�Ў$�l�\P)c���Q㧐F�)�]䬵C�{�sq:��I6<��鍦�5u�׳���\����E9��f��%!���#�n��y��--P���3�P��P�ywH�� ^"/:"
��B�-��Nv` ���rl��(P������u���M�KIש���/�J�Z��W�0�r>����JQ�6�z���E�V�늋��s+)[��{l�KkK�f$ v��K_</1�I� �����:�/N����߁�n�7��_�}��~]����m�}�)%�o�aw�B��3�K���qy'DĨ�������� ���O�6����?U���[{�IQ�cP$�7)�r@rw.HM_Q]��Ugt-�����d۾�,�~u���W�L4R�\T�C��aH��}Ƹh��=���A�l^��4�C#��B�^F��8�e�!�,#AU�罽�� �I�KsA9����y7�/&Ȁ�1=%�꡿��Њ��qmJ�����2�����ڜ���4��8���$
�	����Ke��3��-�����Wɓ6�����q�K��3��ć����1��qW�iZ_�t<9
d��26H6'�4���ؘ�P.50.�Pȏ�����'q8X��X�ύ�����X:
K���]�A����\������ݍYNI����?�RV�Bn.[��v�j�v�TU��7�3�({�����cC�6<�bk��pT���8��J0 ?�hVn�~��&H�u�đ0�	c��K�(ꙣ $���ŀ��B��������~�I�Pu}_ש9Zp0��_�ݯE;��lhlV�������v�hG!�׊)��m��9�g���l���������5�����ݚ:rRPR�qp`I�~�����gQD�G1h�l�a3���F�6D�����./d�D�����BY��ª�a��F@"���� ����>�B˳���#l�������TS�law��B1�娉�c�Ȼ���+��f
2�R]�0�V(�&�`�콴f���9�!��+�~�I�k��RPO��4ח���}C��3�Uf�l�*����]�cl�����ҩ��=�����>��� �l~��E`Z�������G��'�<p��1O�BUS<�`j8cy���h300m�!��ޣT���vG\����̯�1�ԑJ�̴o�Uum�bMu�8��Ǎ��tt�
��8wf�Fx�O���V,���i��璁���$��IM�8ч�:�V�-��o&�z����lP�Z�?o����E�����d�B��@k����:�=>Yh�Ϊ��ڢ�l�o��(��"�0
�C�"�6ReW]��a��YZ�*J�	~w2cݻ8����y���Et~C����X0�(x����8��4`��"z�
���PH�M�CN���U�=��vʮ���Н�	��X�汼�U��7�']���9�af�$Ix�MA��Ҟ�#�P�%m����"�\\(�4-1��"B���n�$�MY���/��sX/  777�=]�[90	��	O��o�'/yE� [Zm����zF�u�C�r����s�T�C!�u��Z6�<����B��~le_$�ϗ��ꝰ�4\��*睾ѓn�`��/r��l�#�p&�1s������l�K�F�@���g���g������f�
}x��	b��QWLR�s��0V�E�����}���]	.�XK�/s>:��\t�)�`ؿ�s�>yX������@}46����l�PF���\��(�.O>����k��o;ŽT���_�
'���8oy�?<������B���L��K���nU%3�=�Is����}Z��B�\f����â�鸸�%�:jZ���ҿ�T�����L�/��܄ϖABy�H��c�� j�c���+�������;�m���<Zo�7x��2����ۋN���`%Eo6\@t*�����bf����;94��������:��})�#ޖ4����	h1�CG�(�L9I:�'2"�E���_SYَ�v�'�U�z��Y��eGOWk�����/��EMMMuI|����X���h�۠�KZ�41���
��u������:H>�� �GS����(ɹ��G���l:�]�#��
&Am�5C����Z�h�����Л���ľҎj���7Xd2�GGj�H�DI�F&�
�=%���T�P����ӧ�Mo2��$�M��(����ߩ�Rx=1_wN
�F�ij.֌�	�oV1y*3��X8)!~����5	�O�o5+�&e!�x�x���r��v8�����ZS#�"���۬�ç2����}���z��L���|c���b����xH�>���IH�sZ�Ľ��
�
� O���� Y��m�OO3������Xz����f��3Ƈ.������^�i�myy�s3�Q�D�
)�4r�m�:E����r���zKW}���wO_	'���r�7.��������z��M��&l�	�������E1~�;<8j'�G$�x'��jqe�CB�
�Q�5𴄺�g%��lx�9&k��)�(����"�%c)n�'3�#���8�pM{�@���7\vT6��tB/���Ek��������;����C��Xw{����
1�*(H�2�ڗ�mؕ�ԣb��nv����F鋒³Q�J����Z�N�<�\D՚WƟ�7�מI�gu�?B�N��i�pu��K����_]_��q6�OS$����qF���fP��P�JK@��`6���d��:��$&f��]?����!��n�n���L�R������� H�4���*��QU"n,��G�B�ڞo��X�����%�����EwS.����!����3���sݮ�S**86�I�B��gK�[�F*�nTH!���nmcs)�v��|��\)��'K�)��/�Wtq�I�5�n������`˭���ڗ�Qᚚ_�+k|��& �S�(=�c��L�����5�C�]o�w�z\��,�����y��/��{��Ξ����(��V�Vrӵ��a@�G�M�J;W��Z��.ټ�lk�J��~��Srs�h��T�A5��h���K�������j���$1qL��>  G�LS�����k��bG���>��h`R�PZ��ԣ{�%^vz�԰R�*@���RI���{0��Z�:�f\��ʋV^��Ǎ�k4X��E��J�i��wZv�N��=�jdʌ{����$K�߸�yuu6I�y�+��G�*N���1C,�_0ыvZ��j��4eyö�O����(�e�I�\r%m����x���D8x����֏���w���bڞ��;��-�`��$t��܇��i�H])}�x[��2Z�!C���}Yd�������撥��sXB����ٲ�KZ_�
j��XY�D�(�Si������Ru��k������(r|�R�=����E%b��WBs�}��G�;�������j�vc�l%/^D%KՄ��RF�y+9X��eB�A��᳧��1�]�-�E�9Iˇ~#-�<8�U���ɔ  �	IO�Ҳ<�CJ�Oҽ�QS#oֹ����WߔwMʗz��A��:��0�� #%R�L��q���u�f%��_W�Ob{�Ij�ɦ�A�����"~ ϔʮ��dcu��r��	磡�=����yv�/���c���q�w�PS�u��JJ���]M��n>���E4{}�0��d�!!�9�8±��G[��Q�!g02���j���WᙜT���/l���K��x�|�=؋"����BAA!\D��#��z�����0Tϊ=ԡ�0�� ���2��jfq��rQ}1٬�(Kv���'� 5���|��������`��+>�Y�������>��'a�E��U��w��6@0�h���eg���ݵ��^��f�\���UȜ/��{������n�$����y�*<�������˝�T��5�����y�&�2���?����«���w���rM�%p2����bY/�Ç�ࡃhEܬ&�j�ݿ����:*��흂���}'\�,�u�>#�(29�x}���s�C���ţc�/�ɣ�P�*d"*��Za�g����{s��e�;9W3�i��~��¶���p44�2���L�M���l��ҡ�7im���j�n��Y����Ǒ��4��Piv��$e9Lݯ�W���vr~�M5�Է݄f��Ԋ�E32F��_.�%Y���r.^�`�[��߬>2��W'�����2�rm;D���%�ms�Q�_���u&��E�3Y��l�&�8�o�p��+���v�� ��Ѳ�2n<�.����(��c4�R3jN�%A�O�]���nώ?{(R�g��|tEa��9bd&����Z���-Ώx���<΂�F,�K-*�"&M�H.:�8 ��_���l���mU�a�@?}.���vt	�$_�2���t��\��ZRv=��VĤGKY�L��F�[���x)�����#��O"S��c����	c�+���а����� �S�k� �!0z�s �pL��~xǠb�{��ѭ��e1쁴��h�t�����N7Zm��J�^�P�r4$���b|�K��0kɎ��v����|8����y8��ߓ��6��A���98�w�(�H��;c�}�f��~l]d��hId�sYZ�+��(�R�3���!�|-��d�A|��{����-�y��>�N�%������޸�ek+�������� �� qR����HL��h
z�-9ͪ�NZ⒐�֪Zj�o���o��,�{���"\�Gm8��r�-��~/�U�Z_~��0u��mŚ������� ������"+� R�M��TQi,3^"W>�*oH��g:�\A��Е�Đ%X�4�oS�gt��)3����d�F���W��⾓V�^t���wk<N����]JGmd����M����������F������ˎ�*�Lӈ����%�Q�㦓s�ܖBס)��2{߲Z`�]��Se� �}��'�ĩ¸!_B�*խ($�C2{��0&ov��Z5ܺ�j�����(�f;swe��^�&�HQaR"�26�v�j�S7���L�i�^���x�딡�A.MR_�O��C����''���W��V`%a�+;9!`.dr֟;q�zK
[r�sw�|-�EN��5�_�7kz�F�+B�*�\MB�|&�4��������S��^�����v�~E
�J��b���9�e%}Q���&��Ҷ��î�L�t����<֟9�e#W�ݑvo���*@@T���7�sτ����/D�X��B$#d-\˲^?~hst���V'T�7�g �}7_�G��ѱg��� ��P3�-m*�8��s1+�vxq�5t�߻X��;�TR�Z��w%^�tO
�ܜ�ſ��+ec�3--A�l���<^wJ���H�2���VVVv�<�((�nn�j�z�KK_�ng�otOd�u�^;��p�-��/�jpH�+��4ѳ����\|��26��Vju��V\��2�,���A	�_@@���*nD� qW�:��������ֹ��D����!yǷ�:���I������>�W�LL������7�6��fޕ4��v;����ÓH�D�9R�,T�eL���v��H����K�M�Fl'�5����Ҧ�t�j�!�M�E�O�񖪊�C'���o_)�_(����&� GJ}?��~:Hq�B�c�� R�*��K�9�K��O�T�D��U?h�xLk&9�v��F��Nn��Υ䟇������0WW[1�FA=�����`�	e�aLnCE�ktl#L�����
s#���oA��Ԃ����/%fL���--π�»��Wi�H59m�.:�E\[畘����'h�`�Rg��L%A����y�u��`g�D�� �*��˝����s��JJ"u�q!TWW��Y=D���1B�FD>2�`�ab��x�����B"X�<�t���j�m
���
����M�66��Q��$�}5��~~Ё�
�����-)��o|��6��٣������:>�����⟇PV��C����"l�$6K�iϰ�} ?숦�׉.>�~[�"�ߧ-I�_W_ϊD�e����證���w_�m��<�W<Jx��N�Fܹ2��y�Y�� )�����\�ޗO ��'�,	Ou3ۣ�;_$f33g��	w�ZD��]��A����uw�U�<l�Ə�j<Z_qyfh����#���Ak^��ַ�i!���m�EsI�V���%!�U��7:�d�k���^��`>�'������/��]H�~�/��Ǩ��	��h����8!��D�u�_������F������or9F�|�?�l�rw\\if��c-�/>�B�r÷�B${5���@��X�d�s;�*����{�AP��St��`��w�@<At��!6�۠��s��{�2��ֹYg����ME)f8N��ǡx�BÈ�a��xmWW�O�����TJF�T�Q�g:R��	�Ζ~��S��_�u��k���L�`�����A�i-w��� 7��R�Gs�7�a�9Q�3�qև�Y�r����{+�ՕV�WU�*�6�3��Ë�<6ฃһ4}&�>��`�Э\�����XǑ��=e\��֙wz}�V��P�G����=\5�R�R�1ق+r�FBӕ?��օ��?���y��D�_\ai6G�3@�.�߄�'Е�6������K�0�=
���d�Y]JA{��X �u��������+8�x/7��H69ȺfO��ե7��@-ϴݟ=�5
|��n6�	�����]CW�i�՚�婺R}"����:#��?��**�M��+G����C �Ƭ�&E��պ<ޥP��6�R���#Mg����iT��ZY�.`-I�Ϳ<�+C��w��A9��JY:�߷sMP�͟����kuC��rff�de���n�m;���e��1��q6��8�P*��V�2UtѴ\S��)p�k�f
�e��7�R�/��󫄣�a`o]� 1d>m�r������*�g����-`��:�q	۠a��q�-��+�ۜ�{?���`����(���*��xz(��v/6�krqw��{zzj=�-�� �
�������r��txThBrD��!D~��#�M���+�trs}��:q�t�� AP�
j{�D�{Ƚ���; ��Ω�ɟ��sq�gbvP�[][[���G�;2�]�δ�Hp8y��f7Et�ڲj8��.FE7#x��~pv6��k�8���Uڛ�Tlg�{�^Ht|<�����?
�g,MO����
�T��j#�F^�:8�眲�-�K����ݯkԈ.l�`�_�Nx�MMM�g��E7�!����2��8̻�m�	��ԩ<��F��0���G��T��ط}��h ���[��c�@�{��N�`W�(0��,+x��*@�lx�*�j�M߀6?S�����m�峤x����ݛk�\��9Y���D�9�w��O��딉QT�z�dddd|BB`C�Or2r��J����o��|�z�!3ׯ�6��n�eI��� ��H��[ B2�Б�K(�Zh"��ܑ�3���S'P��ȸ��a���A>nbM�-ߕ��j�h:��]��m��FHX��O��"g�ˬ�>3�U�hʌ��-��|��G'5ɔ3uh k��%߹��(�zʂ-���Ή�̈?��BΌm�5�Z ��\�P/���b?�
@5��C�ϱ-�
 �� -��-m��kP�ܳ�R�;k�?�Č뗺�M�U�T��+3��B���\ݬ9[6�~Ⲿ�hf�98V��3G���;f־l�����A�7�޻�����H��Udgw�$�V�G�4y��0y'3�O���|��ٹ�f��l��D��ԓ$�'$
q���Be��{Cuj�m��ny��UjO\����X���Wd�4I|"����'��bˠ��K���(�8����w�2��j���$h�P+: 2 �8�Q���������H� V����-��5���X�G�Z��EaM:Ȋ�Uv�tF�O:E:A����6��`f�3wyMA�M�+����t�
�O5~�O�l��<UK�-kV����#6��<5���;��)��1|�s���L��ӵi�f��������õ��Qc"�	^����e�m_��4=ok۲��k�<�^ c`Q��py^v^�0������cc.˪?�2��y��{���#��ׂv6	���b��B9Ģ��U/��v�N�W��-5&�~V�M�����S|;%����l!��T1�����w�2C@KSHp�Bybߛ�$����1����t��b4��a+-�����⪱�7��	�bR�X��EE�Ӳ�N3Oڝ-՜5e��X�*�^��B2^/"�Z���1���h�5ƢtJ��*�;r�(�#��F�`��~�bI.B��, �r���X�J���EE�i�d �w�ǂ��f��)g��p7_n�����߸:��1�?�@'���!&�8���vS�h�۞����n~�p��'B5��
zݑF����?�������0��N�^aX/���_�C�k%����:~<��%L3&�������$ғ��:���ׇ�����~��Dw1�9���\�&O�_��o�mj/�H�֗f�I��l^|i�v�s:M�X��
YK`��Z!�7���;��6l	>9,U�O�&�R	��-�y}9�7�x�E�^�|hϚj�S>�������C����� *;�C���8�f	���zV�(B�����n�5�<�G��H�xa�P��{bT�b����YXP������X���������i�q�ܰ��M�V-�hA�6�H
�cWb����j���lТ��g��w��qk��}�fX��]�� �<;PjP]��j�������T���N�~�z��b���h��!G�+�\ĳ���|�6#�|QH�u���#��ܧ#(��2�~��\�I��v[���@q�Tg�"pz�����UʴV(:�6���V���z3V�C �f.�	݂����o��k��I�����iؤ�ڸqҰqc�Nc��m5�m۶�o��>����̬����`���ꬸ��X�L
�mzq�ԗ��}\�#�ϟ�iQ��~��^7�wEb�H��a��|=#i�A�p'���?Ek�|��� �oZ��@���Bg�7�A���fP�P�����ۯ��$7�	ڞx\\\�)�8�b����Ju�S�U5Ե��_��y"��scy޶[Awm/W�6N&��Z����K[��x������o���x��_��"#�.����:���'��y�������M�Q&U�|�����73��_0�3�)@�,�Y�Jf�jD]��Y�B�)
�d��Gw�-?���]t�&-߇��	k��ENx�������Y���Q���J��ױ�L���yJB%�� �������38��a�3bqd�Mu~�tv�l��j�p\����D֚*)�~T��#�]�6?�7[`sE�u�*=�Đ_�����9�R�-�*�z��Y����be@�K���2��<��y����a�Aw$w�u��Sp��X�A����׼N��B��M�
�\K�� LL�_ ����o��ɉd/��uR���@%�G���F�:���fFmo5���z
<��V ��U���=�"�Kzq*#Vzzܰx���i�o���:P@���ᓍik��G&:f�Ka�7Q9sx����1D�z�Uu��A�̢�jb]]������/  �a5���b��c����'�.~rQB@��r�z���_�.���z�����R������f�~kw��ˬ��B?�asS`���k��o���ӧ��|�j⓵�D�o�&oI\�� !��S3mʓu�C]�T���˞��>[cf6�k�0&Y��L�+5��	$dk:���ԜϘ�c�eLDI&��PƧ�(��4Y��tGf�m�+����y�kH�&0��pvK�l�l��ԍ��v��r�2Cs�a�����"b���լՏ����N}��χ�W��ݕ�=.�/U����ڠ������n��}3*l��y�k�U|޴��Gb�K�s�(�����3���gV���8�z��}_R���'�l��v���U���,�.�����ܱ%�4C���2�ק�t 򃦸�x;+5`�d˓�$���Ԙ6��c�<��;x]�fm#�=�>ܷ��>�3�j�5*ox\�����B�b�L��l����%�	U�0�뼟�Dh�-]l�l���d��:k�ksW�]㎲6�W�1@�K� ��h�����sѝR2"�	�{w��@9O�ˊ2�=/�fTO����/�����p!I4FaԄ��܏'����d�����y� m��.2�~%��uʉu�&s�-	��I�qT�=��\���ҊL�������KǶ�a��#ƛA�e?����B�q(��+�@�x]ݯ���-0��C��2��\�j�b���mئ�b�-I;����#��"��o1ZȺ!� �Za���.���;��DJ:Tc��FP���k�-	'[�~��?��=F���w�}��\���v�\�_��J'��;Ñ����Wr.�Xy��G�ߣ�hg$S��e�ax?�K,|��J�(�x@��]%<`
ܞ5��r.���hy�N;=��vϧ��P��Hi2;�t�m.�g�����q�hN��۾��f���g9�m �<�>�3��D������57?�{�����2�{�)jrr�jy��J_Y�1���0��l_����y��a���ŭâ�YK��������*��No��ٲtV+�L��kNe���<ҥ�~.�5�&�ؗ��F�Yk ��5�&$�B4��%:�~�T�s�O�*��re44[��֙�#�>8�y�e��1��r��� ��1W�`�Aֽ��ih�� x޲��H�Y���@
qĐ{Xq�H��7ϓ0����_~x�c�ܨ������5>@;{�eG}�eO�b5�ݺl����1\�� �r.P���`�/�(�kuL���[����Zt��w����rv�Tkzhi�:i#�A�sv�씠�4�PQ��ɩ�������F�uǹ��&��js����ؾO�!'u�����mΖ�"���ޞ����x�+���#ۿ~$\p����{f1����fVR6ǽdZ[�;_?;�z������'��p��g:ԏ��t��;F���ǻ��_5���6��]s�{��oph�2��
���7a��%D�\��?���}i����Hm����x�03g��q�<��8�<�y��J1�/G�1�ٕcJ�^��������(�!fa�"%��l����T����wC���KT���v��{�Ȑ��K�R��F�d�x|Me���dz���w�.mťŤ�U{��fo����CC�Qk�|MRT,umm�[qN�ʊ��l|���N<��zO���vA7<�:%}קOP�ā�a-��*����56WAq;�{b"�������v�Rt�SQ�l���.y��[��T� ~zfb�a#�-h+9��Z�^P�@커Ƹ��_��2�H�:WR���7) _v��6�><ߟ5�1P!�/����E�(��&[Kr��&}����F*�[}�2��gcs�!��^q���ysv6a�U�)�i2����њ�Q	���o���X�?/��|���N7��?��l�Ean�:����E�RrfL�OVt1�1���=��2�qRc�R��Irc�L�R���b*h���p	��Y��h�M��Ƕ������S�T�Ӧ��N)���NP}�l�R���_��^��

ak^���?ۍ��u��G��G�:��h~�p�����\e�ܦ����ȸ�҂��S&A����e��|�h�S��ނ��&zv���Tb�8��`�ǭ�j*�ϬSȗK�#�C��u��5^E��Qi�~��y[��҇��\:���A�*mk���(
�� ��v���R�Dd��)6Ts�|r�O����m� ċ{����|Z���܇'���NA��:cs���'ȏ���?i�+�3<�o����&�m��?%3�?�!��9�bA�8�^�g��Tv���L�N�D=�7'$��p��:�Ĭ�#''����)P#҅/�h�D�S�ū�m��6�ӱ5C�]������?�����$�#��;����,l�����	�
��L�*|�rY�r���K����=�x�}m5������V�2� --����B�d�Tƻq�]a�J���Ctu{[i�U���č��P�,�����W�FH���a�D�)!����
q˩MY]͆�r�Ӽ����������^�;k|C�sY"g��D�P�u��y��x"7x���1�����l����t�#!I~�L=���Oi��/�ރ���.��v{ �]�������G�N+�9���tr4�.,�y�{��H'�+���K�����Zy?��=�"��Z�5�?���������<q�d��mxU_LD�pm�rk_M��Mο"[O��
w��u"�殁��:3���ځ�v�5i�S���2V�G
JS�]+��cfXu��愙�_hu���K'%�VW�X)�������s|6wg�G�����J1�Բ��(�6��a2T�;�S�������rk��g���'Ɲd�ZX�ё��u�Q�~�IP7�传\�����q�`�&/�9˳����#��zz��`3Ե�Lo9����+�f��_B�u�%��OPQQ�hFz�,��X)����i^�\�*��۷\=?�_|�NL�;YR?<�U�kҝ̖����ofd&q���@��N��%�H�	���'5��˛kV�-��l�{�@�^U�C�l�ѝ�L���'
*�Ё�"d�b-Z�ٕ�-��B��z��t�J�둌�����_WGG���;ӑd�\���%3v��C�B�_��Y2R���|Mr%135�|͗��|]��B5I���'������t������h<�0�z111���mfi)"ۿ��Ϙ�~5'b��ДC�Ԥ��Ē��DW�M���μ��%�U��@ti�J�����|u������D9�x�d���%�mk+i�2��� �8>R�C���_��f����nX)���*!�S�/�͕���w�G�q�(�`�ќ���
��6�oWE�_�����T0��"�=� l��'���t`�+�����N��g쉙@D��M^�(H���w���6��s9�_���p5��P|����EDjhBU�ba�1886v�)��1��B�v2�����s�w��N�I�����XTa��ĩ��?�:3;35��ݿ�14��*�|YM��������I�V�Q˅�x�{wNHL�Q�gn/1�U�I-���u)x�ѿ�h	���n7m� 9P6I��eg�Nx�p�n����5�4+aK��c����s��W:���>?/a�2���jow�I�}�L��Q<(��Į�Kֶ��Xׂ�
����lo��GPҴ���0��î��6D�S��4�o���"���8�0ԯ�ͦjo7��?�5N&@�i����$ۅ�7�=mC��T� )e��#�j]I^w6�25�isib�����5��4����ѓ)+ȁ�F��������y� MM�3��2�淕�J��&���)����AQ���Q�/�M�\��{�Պ~%:�J"'��GItP� �ܒ�aD�`�әz�W�}�TE������f����ծ��êtf �7"M"��ե	�+��1G�/�rf"xCee��g��L�R;u&���k|ڐ�l,OEE����嫙˥��C������̊���Y�μ?y�6'���~�]�kk�����Vhg�?t�[s����׬^�)N�
��Qe݅E�S���ʛ)2� 1~]]�ub@S�����4'Šu��5-��o�P>9��r4vaB���$Qw�!�w�`�	�D�|��r������]ܞaͯNke�q?G�	f�0#2D�S�h���2��W'>=W�e}uU�~�������#�o���C>w��,:M�?D�_�dR@Sr|���/Q�F�q?�bD�fs���������O���(��d�0�z!�MPo�����.�E�^烙�s#(���2#�P8Ի�$��+�'����GW؆Nrdұ=���x���J:'�
.��#�ߟ&5� m1�,x\p��$�9I��o#�������t����m�Lt.39�+���Zo��?N�x9�<���`��
��<wZb����R���6.�5��d:�e��9?����fipY��A�Y���#�]|[D\� ��7ff.:�%�0�'$��G�"��|�|��Jՙ�id]�,��8�6�����a�gv�F����"��-�ґ��f�Q�+�t�%v<k���$�ʉ��&�v}�o襥�X��%��d�ׂɡ���xmk(4���/+�Ε�^����ˡ!��
���u�&�mT��@�w�˛'+WI�<<v�c"B91II;��5Մ��4��כL��KG_���e��������3i���F�`�A��hڷ�iX�l8���������<3��+���y�!����|tOt���9]9�S� ΅dOC�����!uB�з'����T�v�»�6pI�N����i��$o^+�z3��T�����f:&>��GV�kXWV���"�}Z�ު�p���oM)�0���g7n�!�R��.�jv�ӽ�,J���!��"�\�:s�[��+%�v��L��>Z�-Rai�O$Φ���4��%Ք1��.q�)�oʐȷ̧�맪���{�R�CWz�
ֻW�"� 4�TsL�9�����[1���7�o���)���D�rtxٜ�%�(���z=�E���c��"_خ�#c�4B����D)ݣ�\���tNӿ�.$��Ԑn�o���4�~�݉	E��In�v���6-�j�#���KK�
����
r�1���|*���Y2�����B��-��� �."�ے�I�SNYI���m%�������1jZ������m��z���w���0$�!{7ԸB�`L��Z�F$���>��q���ts�Rz�����~<���,�7����zB<�҇<�Ѿ�X�@)��
���5��ۋ�����9��q��#�^�Tq�����?2E/rσ�e��V FzG� ٝ�4��� �;�a$,7�@4� ��'WC��{�%��ru���i�8�@������ 𷨊�ܜ���2�,3�Q��Nr��|�7g�o9h
��ؽ�~ߺ��u�_��(Ak)����P����!^V��:5��yAT1'���&&&�rj}8LZa��Ծ�%F�ڲ�\�+-SC;��($mɊ|�_�c}��\�^i�*b��������Z��#"H�R�|m��Y����	�۵����3s��L�h���yyLn9X�]����EGE�����U>"���Ha�Os�|G�urڂ�F�K�Rt�(�7���3�I�k�̖���ŝ���0�͜����s�Ū2Ds���F���_����I��xs�p��h�4����oM�Bv�HnY�g�,�^f�d#U����gtW�rh�K��@���:�Q0�S,W��l%�g̛�_mB�:Tj���F55JW�٫̥���B�����td��Ib���\��y�s����z�Ũam�c�[#r�`���_Ψ|&���0��Q0AN;�)�%w1���I�	U� ����o���YX\�H1�"��xdj��۰/u��|��ܿ��Ĵ���p*��#P0K�0ANr�5@�χ.. ��/���I�g�3�##���c�%���:T�R.]T3c�ͪ�bb�bc	�������3�W�^��[Ӳr�s}"q�-����S�I#hh+Tq�]&]�i�7D� T����H=�NM�0��X�����%o]Q���TM*�x%��-�I-�l$��ަ�H���Tohh�����Mb��?��m�݆�c��.�f)#c9�X���Τ�9C��P��͍ا��/���I��w9���ޱ��C$G���Ώ�;~�.�������P>�ɋq���D�׽ѡ����p'�:[��u�yV�U�74�f�Y[���ۓ@<]p3d+�-��C�t\�Z
��%�j��t�G���%M~P1�����P���SKI�j�lw`��̘�`�TXxfvv[I��8ue��-w6gkYu!��l�R�r�xd�3����cvb�ik���p۵iQ x�:XW��*�L�To��3��d6�[�����N(�P�n:Sm12�~�2*>������V=���,&��33�e�R4*��3"��`2���t,,·t��E� ���������#�����p�o�P�������ggg�'"�����%�,6���<���zj/���0[)��o�(�����r]]ae��/cP��R2<�.=�^���D)�m%����%�9\V�� !&9= 'k�m�� W��á���O����x�~�Y����C(/�.),�c�Ú��"��m�f�ƴ�U���.��V�I�wm϶l�	�%5D�|b�xa4��H�:����®�]�3�(�Té4������;de�$� Д���m͖�	�z�[�}
����Ӟ����"[j�����с�ךĀD*��$^�N�L�h2�*4�-x�8�?��P��SQ��K/��5)���T	��ތ5��eS�Z���� �����Q��VJwQɮ����&�t~����k�!��)}�ar)i��שȬ2y2 �^�ie,�T�[��Xu��.���P�_횂g�hM��lE- ����/����%nKM�򢂒<�O�6J d���ߌ@&���`���>l���(ܫ*155k�%켕��5�N�a�=M�0~�!��G��/���hMW��'����ո��iR�Ww<[��.1�{h{BP)�@{�Αg��C5��܇��d� ��n�=J��t��F8�9C��u&�臐o@rr���xQ�̲��?�9�_�VﵕFŰPPP	.ư際�۹>W�ω�o�ֆ�683��:1;19�;��k���Ғ���h���BL�*]��[:_Xi�ഽ��#`��#0�����9}=9����B��%��5��T�l�F�ʶ��۲nnk� 7�8#D� )yP��.ڙH��e&�;�[��QvN�U���{ȋ(�w��C�Ep�R�x�-�M��qf)�vZ#n�@����vw���#ڋ�m\~�F��Q+�����3&ymn�JQp������x~Ѡ�����f����Y�($ߧB��1����6SOf��٪�{T�b���#z�vLO~F�8ؠ�ٗ�)�W���"� �t�e����ɾ-/?\��U���=<,.�b�m�xC"�a@��vrr�(������:��iV��?�ol\Z����&��Ge�wπ���"��p�d�<@�bU]N.J���i��=����ۀB�N[w�6bM��7*�L��s\��ʺ��aOh7ÞMk뗆�k����R"���WZ1IJA^NZ��O�S|!�}����9ЇI�N��3�����['���Jj��u���Ĳ��b|��׿��a'�?��,���=Y
�2jD7�Wt���td�)?���=��4��Ņ�{Zg�$��]��W�S`/Su������v��}���E��m�C���ݏVw�]�05�	�`Ɂ��n�,�������H��5��ݒP��1��_�8��'
�,Y
�JEq+TF�L��݌uR����º��#-�mQD�Y��	sW�C�E���<�$�:iZ�Y����Tĝ���i��
r���x�	y���F0��ik7�U�!�	�ޟ!qpp��''%%ua���?ř�re��7�A���@��?�\��c����h�TO��h�]�w6�A1����%h~�k^F"u������v����>�P���U���b����}Nw�V�=�g2�����
�U� r���0e��,G�� �Y����kD1�U�Z��+*<��#������I���	����Fɣs�Wt7�u�P�Y:���]��(���������-��"ā�f@�?��}S�x�𧋜���/������E8�$ܬ�*�&�,+˧��^P�$Oy���mI8�g�?s����)y��B?��j~����K�>�{+%�"?C��Y�
SY ;�/�A���矋k�S�ϟ���)?O'n�����AU�#�I@e0E=s:>����d"q]�hk6=����(<B	�ab�o*��HPإ�����yIk��pTr<l�e�Η�S�OF��c���񳔣�L�5a��v !�Ƕ��N;ft#�b��Z����%%z����ۗ6W~j�~;;� Z��TxS9�H��g*�r�)�Ӕ�b��՜y�#��L	0b������9;8D��ɪ�#��)�m賨�%sSɀ�-��c�J���JLL�BXjz���y	U���gڱh�1�#59�&�c�T;:&��X�X���.AHy�PR"�҅䘒/y#l�N�n�}�N�p�����4�Z���J`��~vS�����O�r���A�o�L��G�>��^9����!;�4zH�%�|@x����|}����.����(�� 6�FE� 8|l�� ��po�_Z�g�0���VX)��n]���C��97�XĢ��kʍ�{��s|�Hm��%���XOF,'��������G�9����kl�X��E����ݮ����)nb7$a#M���wpaD���}�0e��;ڢ���֎����^h�&�Ϋ�2��夬�Ɖ�g�m#q���= �%[��C��0R q�)���)��-��1�2�6��p�i�U(��j^�ҋ��]�vp�7���W�4�C$i+M�EjM�e�^�p8?�#�����N�w��h��C w������x(�jD�ק�i��O�)*l�4�j�h��;yn;q;οO{?g�cN�F�.�Q�[<w��NVn8�;G�H�%�'�.��S��nc%6D�E�#�"B��k�IV����\�Q�v^__WYova�1��_����88�&��:����D�Zn��^��-����L�5O4�{§�����>��t��G���?i
;A>��a�����W�~�^.90� �������	Փ��jY�9��x���O��i��jN����7|dㇵ��ɬ05E���ն��۞�m���
�=2�����70R���J3cNf���k���#5a^�)e�X���U%��*��M��>��ܓaT:�`bѝ�(�W.�DJȅT Yi��a�V�ݐ+����Ͷ�1L���򽦈8����̜��>��ݝ���˚����Ռ���g
(�<Sr�}���0�$'d��3VՇJ��V�: Z�Mt��kqM�Kݞ���핥O^��OӲ?ϳ�u���t���U�NookR���qp��Z\�|1NV��3i}�Ɨ�;�N$�����+�����[����3�J�U�^�].�.W�m׵��Ǧ���g�,��b��q�2;�w&�?�?�_4�@oF��L�H�ь���6>+h���R��HǊ�ŮLe��e�ڧ�������`�m����8���m�	c�U��U�����?'2��C{��vؽ���{�p��b��sA�Ƿ
�.����B�oMUڭ����`����C?�D�O�ge�KĘ�cQ��}������.��n���x�U�ʦc��\��1�y�G�"�}����+�3�u��̂\_�	=���S2�n�1�-�E���^?8���9�� ��ꠡ-��"�h�#�W���p��P:�xZT%���$B^^�Ĝe����i����!m8^P���C���;�������wӸ<J�b|n~էWFE�V9Nk�tf�w�����s9n���$�XXX�~����Itε�_r�;���E�:hs{��u����{����
���[��,��:�dk8���7<�yR���UAh�C�&R�fpG�kj����R�d�)� $9t��!�$�{o�ާ'q�3��m�hBE����ɂzjHצG�@��^�c�]��7A�ݺ�ߗ�5%sd�o�}�~ȿ�?@A� ��yZ~�-�i��Sb�2P��@1:�$ /Ͼ|e����v�
�{r���y�Y�L:�{{�"Ķ��Ҿ�N��y�� ��"�|��i% �'����n�B���"�~� @��]L����c��f��k깸45�_6Ɔ��M8ԙ��~�ׯI���ϖ�X���&��|��h O�5�w%�I�wHUĆ
ȋj
u�/�z�U�KWqq����d{W��QaΥI���OT�=��E�pI<�^���,�-Ʊzzچ52�!;�.��jHI!����&o��]\�B�&jJѮw����3���@��Z����S�=����$6���Z/>@�_�j���T.`>�4� $gI��u�l~`m���\/̜r��)�Y��\]IF��&T��NM^��Dѻ4�K,���;1>�B���M#/w�U��_K@s	Ê��1��шTā�1���%��8���P8��\(�&s�_� ts*��2#��ZJ,�/�������q�3�����1����ژ�#T���x�����15yzr�74���Ę��6@)�4-��/]* �"HD�<�J�	Aɞ��z�[������x�_���(��;�)��C���ߤd��h��k;x��'�R��q�l����O/CC�;{	JG�v_d��X�v+����3���8��̜��k������>cv��!���[;T�A�H���3�cZE��ܸ�?s)++�~5D����ص�NN�.��iP�
�@.��oo��:,Q*Q�Y�Z(E�B���䄋�O���3_�-&���ƻ�T]�K�{(��
B;o��P��ֹ�g؁��Āi�8=E�����/HO/����r1�RgmW��/���ȃ�a/ߝB
J#rrm˶�N 3�����c�W.��T��m�w�r����H!��XT~#Q	a\��� ��qa���c�j8��WS�q�LZ������׋y��\F&��G��:���I{��p��r!�_x��������kp��/;t�rc|�jpD��ťJ�W�C����\��>���^7�>ʊ��������eύ$%�y`l&�� ���!1�P�)9��3��i0�B�Ʊm�86m[3sY�!P�l�%}����ظ�M�l��~��>�Y���	#��]��?qs�sss?���_��0�[����]���Lp�|�b���rK��4���Z_'q�;A# ܽ~��C��Q�����z��P8��#���&W4�u����i��MIM�ww�$���H%%�b���%����;����Ơ�5�Ȱ��y�g�g���^��2踈܈H�������2������*��z���.��-�)�sW�����˻/���B"*-�do�d���|�[�^���� ^�}$髼�;��t "��ߣ���������ô��)�ڞ����rK�h�=O���XJl�z�ll:�PS*W]P�/,���2 n��s�hWs�Y�%��w���V�͡յRj2""�^��6Ի7�AR���*Ftf&uNvM�����6vvfv ���Ĵ��$�'~����i�Tџ�'��6��t[֍Vyd^����=�e�B��0wg��4��t�wJ::�"��$�K�ۿY�6AYsj4XC\^^N�΂��*����^h���<��6����J�A�T��y������VVad��&�>��}KJ���T�M;��X��~ ���oo�|7[�//�*Kv���U�����0���ט�J*$++�r�O�9i�pZ���2�؃�z���Zk���F�yHl�J ��b$~mϺ=Ah��  ���xt1?gwF���hA���ŏB��0�̆#����:�O�_��z�p*cm�4�v��M)�����
��H d~ ��9�[��p�[hm��S�[@��G�65?��2�㇄�7q������6� ��W�R����F���[��eb�=C��84���8�z�����_~C��q� ��tH}s4���h�M�"�COv������IOO~��!`$�񮁡��uqu��}�n/�HR�}�LZ��r��J��q�sb�#<���F�A+8����+�����7vwg�Y��t�n� �ֆ8O|�Fy�_�*���;^��AFF~ �߾y�Y �1���+�R�vb �ԒiG�h��F:�FS��D�^?qr��Y���&~5���hv�T� �t��>|�\���ox��>��@@Gp�y�����W�VARˤvt�@UO���č�����̗9}81?/f`������c��091�2��*�%ס�"��@n3����A�|2~�Z�)X�L��iv�t`k�G��V,�W��� ��tV���� ��è��<��.\C��%�v�s��|��iW��G�)�Q�H����W�TJ���C�Ĥ��@|=��?}���hf��:�� #Uq1�u�.�����&�!�X�WX�64L�:��v�d|��:� y#~w�rr�V��������z����h24hö�A�?y����"��-l%121��͕v��6O��s�LBUUU�Wi'���T��ȯ9Az�elhCG'��x�\�^���.�Q ���.A�t�s�}q:�@���ޞ�?����8�"�
�R�_�*C�����Xm�qI�1���p|1H��)�����b��0��G`�M^��p�����ब���4��e���F�}݋����Z���H�z�M�l��Dl�664lT��wOd	m��!/�3����묷ypz�8�����C�SA����}�?����c����y �Dn�������<�P�";Ln-[��nt���~�D �����n>'XY]�2��A��&��j���~��O���v�
9q�����-OJJ*,6]Z�Y	�\�@iE{.��~�b���>���P �z"�g.���Sұ��)���ۦh===\��A  Յ1=_oU��􌍃^��}Es6�+����=�!����l�hJ^�

FG�	��X��k� r����]]�������>>>���*Բ�=���U ���$5x<����|5"���E�<���c��J���"�xrs)�<���U�����yh�r�0�e�G�ۛ���";�zC����?�&��3Ȃ�
 �s�����&M"/���g(Tz��k������������G�
a��}��3�$����v�t���F1߅6P4���\Y"�S��B��?4��˸����uM@�, A�M��	�;G_G�ʏpp��"����jq盝���׈����y|���D#Xrr2�0 �̺D�p}�l���	������c�H�������J���� F��XO� �P 2�m�7���-��n!�`��i�{�F%ZDĖ�ͨ���Cqm|u�AR*·��rr��4���.ӰU77�Uۄ����|��8q s;�n���y��M�Z�}��|�����z��l���۩������,JQQ�j�)��mOū��\8h"eb���	7�).5�̂���1K5�����AHLqqq���:Vn>�A���~pt�5[��Z�-���o��?Q���&#�|u}�e���ge���� 2V�y{}�kdt�Dvv��
�ONN2sr|� ��n#� ��3Ǯ���d����Y�ٌ���]Ê⇣�
#�y��V����:|='Q��S�����*�u�ܼ���}}}���p���߀��D"�9٧�' �i!!!A�_�~-��q��(-�?8>�Ex�'#����,���<G�B���F�h?�h�6�@X&6��|��))aKKF�e6�&s��:�!�j�ʵZC�Z]k]�֫��BO��Ɂq�Gijj����r���Bg�ݫ]���NJJ�\Z��� 4J	� Ձ��qoR��]�� D���NM��Ó~c�j ��<l�=��2��iv���T�@�(-�B���`��Ô��6���L��;}a�)��y��h ���F��--�#�l��D14�����a�������8�-���$2Ci}�`�r�4臌L@��uVJ�@9���M������rƱ����=������!)�J�Fg�P���J���ـ���ϟ?�E��&�onNA�Й��@D+�<����*(����tsc#� ��5�����Am�|����4{?'7w��*��d�Ab����f�?ț��Lg ����̂���~��=��W�]}��� ��7ce�;�Z��� �ȠY�|y�I�k��/S���Xf��=��K%p�֏^ߡ;t�Tz�����U:���Bz���:���1�?u+�]۴>��e�����f�SW�>�����
���#A��������N۝� �XY1����A+�,�P�٦�=~��Se###=mk/s+��\ISq�lf]<�!������KYsg�S8��  ����������	#�������"�i�����$S� K\B_��Q'� �v���zg������tZ�OR�}��I������
; 1��O1���ds0A�{
�+(��dЍ�M`󏈈=�ⱕn��=���
Ӱ�C)�Z˾[o�|����_�5�\o'�������Jߧ����,x��2�*`�+@ $�@�K����"\
P>P��S���Q^/��ڡHuPBJ�Р��
���hap�^?$�Q�%�_��R��e��"�|�t���Y�_�"~��6E��a��ݲUPD��#�M@���Q����h4O��8�c�eu$}5�SV������s>y��f��ëz���7y��d-���[�`�ml1��W�s���Թ�%�z�����*�Y�����؎��D�. �u�T���3�� ���Ay啘i�@pڜ���
�c�����n���e�l�X��\�dee%~��KQX�5���*|j��i+�)��vj���w~���M\6SL �m�V� ���: �Bq�� �.��SɼJ�W��g*�ԏ��j�H�"�,)���^W�����lɆ5��s�G������Q���掁���a�v� ���Y"qwP�&d�0t`�	[V"M�J���h*Wu0�hUMM�� >>M��ͅ<古�� 3�F=�.fA�曒�v�!׍��[7!�����[�����M���N�?�i6��7kR�6��A�T#���&����ӽ�=3ihj.�V˫����}�]*L��/�]0�H�'�
�Z���\mr8Xm���c7��ζ5��`���'�b0���
��_c�'42 Y�!�7� ��D���}TF2��3��3`}��Q�b����M���/ =� �
�J
U���?��"2(�#.>~@Z�h	
	�B������Eav����i�i�,f��0�νu�g$m�W���k�JUz@)���94g=�w��v��8�֦8���7m\ �[�^�J@���:.�+k_��8��T���"����+����M�.^ ۝RU�_�1��%�o �V�؛����-ѩ�o r�o��������`��~U��	`d,"��-��J�'4���[,��խL��F���E�B��i2bBBP2�p N���t$ *Èx��#�ȹk�z������
�1@�J�h?u��N���a}ӵ��b`V6J�[�(��}�H���n��dĀ4'x�	}co��3ȥdC�w+�[
ff4666��鉉J��B(��$��fgg���c�
 upq}k�N���8��10(ӧ�Ɛp�cY�����Sf9�#��H�)�ը&D,`z8ȉ�^0��H���z�*��k��-�HH��4"�tKJ�tHI���� ��)Hw7�����y������V�p��k�5��k�����}�H��:@�Օ�`�W�fgg�>O�T�� ��1[eնv��ya��[3��������!�_�{�W�E������S�'(��WR� S�<u���p�e@Y����1�}�ω�L	�jzzĨ��⋁�^�'����^#��*����{b����bx�3���s����>-bzZ�!���/���"���J�Pd0-��m����aO"�ߧk?����Ag/	}�R�6h�*:�	�}i�P�,+�ҹ���D _�JK9D���ggi��	j얈��c���,6���zU;�۠�nL���p��[���Yh��s�MÖ�|�&se`��텘�½� �+ȼ�IJ�$=8?o���ڛ0;���O��.!Whњڋ�=�HH|�q��4�ORX��U��Z.+�D��_ܯOrFS�''�¹"���JJI�pr����	� ��AH��2K�
z�?����b�Bn.Zh}v~~hG0���F����|]6 q�8��f�ی���߿_ �V��!7*���%@���!��z^$�U�H�m�12�Z����yi�̷�����]����˄�kEQ��4��/R9������##�W����$d�����L�[��ru���ʪZn���<t�1ib�Ƹ�O>B2''��P���ʔڱZ���ӭ0^��t����K(�]�������/e�F{G k*u(sp���3o"##��^�~�e��u{�ggn�
��aC��p����2��d^� P�J���7� �+^�<�(�<���I�7X��<2l	��� ZMd?5_���&u�o����~�Ҷ�z�� ��i��\�!�6�_���:!��� �U�|U�e���̤����̷�]�'�; �v�p�b������� ��2�򝀏�UJ�q�%�'lK��������z�֒B�����ut٠b�1#��Q����']��`�����@����ӎ���AFA	_|�=l���5CUg"&G.	�UfB fHx�����WUU��_��K �o� Hf�	�|�����d(


J���.?W�`����ҒLX�+�_��ߩ��S�љ{�k?56���sa���,F���;�@���e�g*a~�����R�����>�"V�.�%q�WO����/6.�A�*""�# ��0'���� J���# {���v��gVV �_|!F`ZQ �N�{@�d�4H�$:����%�xG�&�j�i>JcR���W��)܄Yc��:-��>$��5Y��(���MJ�*�o4��J�:�� ������t�N�'K�ؐB�K���*������ �?�tv���I�-���7.cN���uB��(3��V�0B/���N��X0�魧�=x B���q���8۟���`�C����R?E��շ����������>V���d��v�����_M����e�a��]�p ,!�צ��o4�/��J�'&##�|���e6���2g@� ��H屟��7��[�q�nk{}&X��,-  J�q�a�+
�]���-C�TJ��h�O�'&���P`������C��?"F��FE�)�k��W���m����1�Z����1xw�28^�i_�I�|���ɨ_�w�J�,Ǚ^���v����������jy��f;#H_�_~����!�/-z� ����X+��ڪ���hi�z��GZ�&�&�v�������7�P�\�W�������dU��I2n�	���%:nR2e�o���j��'�ڛ��2�D���=2M���M��ļ��~u���N�G@ƄQ�_�p�X"`�>�:�;�� IB f}c�y�A���;?�\p�?M RJ��i���}�u��<���"����
��3�/�쬭1���k��W�|?���q����_���3���7�����dNr�����TLF�����r��|�����S%=�'����/e-%����<v ��Yzd`x�>1z�	����$hXT|Avjj�/uEE���%�ʹ6 ` ��)_�{�.k��/l/��<��6 a8dda "
���������������4�!~@�� ���x�/m]a����-���KС:�%���wvh���G�j_n��=��{�kD�$"�ku���Vc���-#�5��r��RT��&� ����̋&�bX��i��o$�`3�EB���)�!8	������Sޭ䞴#ޓ��:��JmY5�ϝ��۷/.��٭�f(�T��׎�/��TUUC(my���|/}N���!���e��c�?�������btTrjr>�Γ�?����@�)�8�?^�BDA�O�D_6�N8 �+�9rY�v���� ���W�^�;j#V��D'���$�.�) ����y�	�0086�3i/L�am�l�8�vDD� ¼y����O�����g�5TY_?pTb|'�󬁿@c�ޛj���Td��ӹt����t��R28d+�e!J���A:�}D&f�v(4 ���,;��Yͨ ����{��3;���� Ú�@j�jW8��a�������E)�M�Pp]]]�F�+��n������k6o2�t ��d/saWJ�X	��I�}귄E6���	3�t����.h'oa#8FJFF`Q�q�W_����𻃣�=��V�����>��?Y��`�;-����ٶ��7��M�7t	��qiiQj���\F��
)������S(i�k�k6Q�b��\�h@��;B0�����L������Q��-��a20V��]����؇��M[U���0h>��o��l[Xx
 �0�WIV�2f��1tY�߀����ק������T�W��;L�vs0�ͨ\;����P*���ךz��g�o�]���ϵ|�%��=�-kkk}��jf1�%˖�̆(a��R�c��]ك0I�Ŗ/� �<Ӯ}Ľ�q���O #(��lhj�c ˠ�1�KS��5#)�����Hb���*�cP	�~#;3Z\1@���z8�DPHɟ�����E�p��b��%2$oOOO���z��D�L%x�����4~e^�SV��8�4a��]�4��Жm:����Ʊ�an��C����J��R029��~2�T�1Sa�-j��}	dvؗ���� z��FwG|}��<�	̕o�Y�NJ�G�Ӓ���s&��PFgKGC<:뷎��4�Z䵺�P�H�0J8?��I&�|h}���k\���(e����p/�ܖ m�̒
o�:]Y_�:�6��`�Tۨt4��`2O�f`���6�&эeW!��WPN��C��`�Щz��
�5V�[|��c�\��!$Y����u��;���!.u ����o9(��L@��1	��QO!�a`7_K�?��	���Ob�^��R��fH*�v�++��Ý��lU���=������6�㐳lg���ZF�m����}A�����ۃ����ͽx�t����Q|<=��nJ�;�_���U��i���H�E� ���p,m���:�q���G)���M#g�}��������η�\}��-/�p)�Q��4���B"ۦ� ���9)T�@�Ʒ��pB�ǡE��&�#���sZ�'�D]����һ�ų�V��V�KS��:Uj�ֈT	�p��p?�y�"���Q̊�����L����5q����(t�c�kjj$���III�&&� `�UWR�3�2�i��*�~�0� �s'����D@ȱʿ���fPN�r�`;_��s�(�؂��D�����~���c
8m�2l������N�����B��)o)�,kLd &��k�`V��,6�wE�YO���|�w�:���E�*�/n�`�<Y�ٵ+Q�4h�x'���P�_���#�YY��dܨ��T�_i$ ãZ����r<Y�ZH�P���`�r��R3ٯ���w|
��_�D��ө\�g�E&''��ޕ�z�ﰎ���4R�lŪS��r��}���d��T�T^^�=YLe��l��2C���,V���}nN'��%+�|geTT��xp6\<<ڊҟ?遝��'�h���vc����#�����|$��TtPv��Qm�0{r9U�i�ŔN52?Raoȷ �I�X�{��+�^��e�h*���˗J���nB#2�4�u��o<�,-х��3���=�o��5T�%we��s��o�y#��R�>�=����uhU� �˕$��*����bc�Χ��<�v�@Mh���QEJ�+**����q��=/���jQQh$�DS��T��+Y,�.wG�kV��>+������@������W=A��Sɇ�"K++rk3N�:������M�Dd�0���/N)�������KI�.*���'����w�n�RWW��K>�� :�(�c{$����z ���%�hJa� �L��7��K@�@!�ˈ������΋f�tk���QڒkU��Ĥmj��v���u�L� ���a��jXZl��Ţ+5�^}�8\��
'���~4?>x��b"C}�3���g&] �E���)Ҫ��8�!����� �(�H�ٟ�@�8(0	�`�z�(�	e�ѭw���� R*� \��j�p�L�����'���y�K�ep�7��Ćn�DhEn�Ӷ|�J�w�9����0Z`آw��X�
�#������4�q�-��YBB����h�撜=��X����f�\��9��:�G0?@�����i�<��Np���c{GG���N��J��^�җWUI��T����-E��1�����F�*� ��Q��3�^�w���w(0�B��x_�ڒ�p�W�q��E;��J���]:?]����H]�����^�.S���npp�+��^d�����Lq� �n[
?I�n�i1
\�I��}8�X-'���h�N�D��囐����"(x]]]ta�bb(|�*������[|��Z$�W�/�����:Zm�^�W��L���y�2��Z����nE��L�l����O����4e�v��42�����;Rn,}ww:��硑����7)�*@��ֱ��o�t�M�l��4	��X�*-�ZW�a0��%��s72*�E����<�h�\��&
6
���ǆ<����ߗTЅQ e�����PmB{����Ĩ���*F_�c#�������@yf�[���R��1Kg�z�wB�V2�x�Icc#tT����۰�$��������G��@L!�J��eJ�Ϸo�����O���%%}��^��о���2E���@yI�K�y�.R|b�P.��c~~>t�8�^#���#��$�O�R(e�m���7�"�;m��|�X�O��ð�̟���`�TD���Ąf�9��TAF�[[[�0�����Tw����dX����wu��#Yy{����XX<�M@W`��4b ����0�R�g����l����wc���8k>Nȧ�~�2tpWHW�xJ3լ��[��p��e-s/�}�_͋܊5�E��������JGGW^h03~:8P+���3��}�&<!0��}o?�c�<0��}<|�aD��F5##������y&
؉d�dO��qO?�Cs���L	<F�3?���

�њ::�'�}W`Ԓ]��W:�{��D-�DLdde��
� s��B�#���Fjj� ��,O���M@P�*�����_deg��$��U��<�9XS��+!����.������m��ʧX���<C���[J�^��ߒ���>�D�W"��8���s����pF���&M��xn�U��r1߿���7��O Ôh~����78\l� ZVV6^ Q�I����n@��������ʇ`'9q��M�P��|^�Lb����(iȟ�jRf3co`��E-ţ�&%$�<��Vd����+�ɋ
�����]�UR)UVm�Dv�9�H�$�D�&����y�α�6��oQiV9^����f��<t�� �d��AP�9�Fx��6��m �$k�҄1@����I���������g69^��&�� Q��|��KDcF��|v���Ӱ��tgX@霯�vK��s5���MLh��P��$���FᎴ*L3�bl9�qjh�8�y�|�|}bªרYGM�;����H����h7�@`jjk���S�������,40�nB2����RI0+������@^��`�ݵ�y؄���U7�z"�\��J [@�CE��g���u�MPk��.V��1|"O���"���7Y�����s�茶���@��𼬗g�<�����7���mUPsa��,����Ӊ��A"c��e���>��@�M���:�NE;%��Ab�Ss~�BK���;YY�΃B}��:.4� �����V?��
V�Q���I���-f�z�����Y��u�K%(S�'pQ�|��LP��}�����m���=�n�`�4 ?һ�M���A�K9qܔ���/�0:ɿǇ����[|���~(G@i��_�i�>;sZ̫���;�,m�Fmİ�s^�nIa��ڿ�;h��$�y�l�6�k�?sY��e��]?��W���x+�r��u ϫ�as�B+B�0��rb�q.5chDE�1�--6��x�P�e���=?����-�CB��t�=��;;ˎ���^RaS1�l�Ժ��46
}�g�q$�˞x�b�,��,��T;�ꐝKg��TK-��'Ж;�Mʰ��f�Rf&��)		��Ȼ?]���������7��YT���{˒��rxff����}z�YȂ��C�&�5�0��8�������2P؇ ł?�D���ǆZ��%��G�i�h��a�^j~
㴞愖�o/�ǎz�5@����u���t�Ki)GD$y.���Sg��w(4����Da�^� �H��*��ڕoK�3�{F��ۿ-&S�uysP_D�\"յa�Y�R{�N]�h�̞����I�ηD�����6�r�i=��ÉW���K`�����Ή��9��q�j�X-ޚ�=�v���=�����u�H_]1.(�ϝ�y�G�\���Q�):!�!�I�$`�R�ZLtc�qr����/������V�cb1̤�s��v>��P��<F�0��������}G\�8�)��YuxD��O�=48�@�J�]N�G!8��:g鳴�,�[�3�s�7���b���D�Kv���h��k=���7���kٖ� h�r?��Vן>}
��#��h�Zp,O ��%� I__�|V8*�����:0{񝓋�/5�) �@�&�<6R<�/ (6'!��'2�`��<�2pZ���z13��;#�g�U",?i�w����R�`��`$n��4�̲NKcf�@�>??'	�/���������������TQ���@�;q�p�~� �tz��=GY.�RF@@(����#X�ːLjmd���5���-��NĆ'�VD�� �c��s������V;Z�D�#����� � E7��_|Z9 ��[|Z��c�5J�	�r���2�v�-�"�I�����C�F�χ`�'�p���E�0�(��:G��j(Y��>Z	���o1Qɇ�;�%��\�����Q�.�1GEm�i b���[��&vǶ6.��N��)�5�Z�s��7-e�,2S����H�N����7a���nh�o�����NPG3�s����pw��\v�B�VSO�pڤ��D�N�O���hY	@����wj%ɹ���� ��>�]���������J��W��By��H���0�<F4q�B��g��B�� G��΅σA���x���qf>�ۤ�x	���hH�������G��	sv�G�g����e����l4����묹~�yyy�G��ڒv���6�4���$&��I�rp`�}������@HI�Λ)�=+���@��O&�O�E� #�*�z �'�p!�c
��ց��Wb��M��;z?1�2��-��J�9�3�����L�ul�M�Ϲcba��z�1������{�x?�]nBiۼ�v?����u��b���X*K###5[�22Ĭ�5:#cc\

L���1�����3fR5�&���~�O{���*mF��yX����d��Д���b��Y��{���{F���ў�<[�XT������{W9�\e�v���F�������2M��'��$k�M�^�l�DfQ���`��Z�=�	x��@��T�Ř�Ȏ���^�b��?�X�t���1}����||��m����=���^y�Tng� Nzt��·�XM�rA�|�^�e핃��׹~���L �Cʼ��3z���ܒ`��;��@ 
m4�����/��ta� �ʁ�	쾴\���@�y3����L�?0����m ��̕:Hj���5[���G�������W��5vx���=���_sVY�Z妖�Auϥ��~yu��|XQ��n�9ꔝ��2U N���ޞ����-L�����·����A�{Q::��>��IL�%������kݑ���/�n�de&�O-�a;"��l��L�?�0������%����7>��@�uUO@�9��dQ/j�xFt���1�P��d=T�����U��HQW�G���#����O_A���xM�_����.K�1^�L;�sE@�-�� ���Hb�	7{�)���Y	3�:�����q+j��\�@IW7i:jj��b���.�)l�'� P����+�x-�=�xE-{<	�@g8�r33��[C�(0�g�x4�rى�uŀ0Q��bbaI�l][[#����r�Kth����4��ta;�ȣ.b}J+ �����"�_�Ke�����l�0���$��-�r�xt�K��π�t��'a��vD���:-�K����ם��P������0b�i k�횯7M��^E��<�4#~,�Z�]:�j1lٿ��A��Uɕ7���3� U��x􆠠P�����o/L�:�}�]U�H���� ��}�x&66���@LB/U�����N65Wi7m����OKK���KS�o�l4��鈺���[uu�0�}�S�%��!�G
���,��T��F�u����J��ʗ<�@I��6�>����b?:Tz�h��Ʉƾ������ծpTTT�H�3 ���y'��L��)}���E��NK�|cRRXNu��b�NÊ@^_,@�(���4*�89q����?c[ɭ�#P��V�Ee6��i�nʻ2�)�i�J���SȭI:5s4�N��a�V���6U���L�]T�?	c��=��kv?ݔ�;��u
�z)�W�W�~��{5���Ӥ����ч%��"�{��Y�=���HL1'�@u(�.��E�߽{R��N��)2�JXtO���8��G���@�-..�v�* �MWYCZz�CUU���qT�FzzD}�{��O˭p�C���D��n��M#�������l��!�<��&""��7�W��j���JB���KH�7ee��q��9��I˼K+�H�w��Ӌ��*�u./�Ԅ���KJJ̿���M-��nj�psyM'R��|,-:�җ��N<�G����8+[[�7��p��|�!�'F�F4��CXA3�P�'888�z����ʪ�|J�^OPt%$��Mw�*�o1/�Ǘ]C�-�!�x�.�u<�������g��w1;�Q��1��N3����k\񑕽��@F@O�b�Qqs�o���m0eb�i�p44L��K+�����Q*S�R��g����'vpQWGh)<�[��Q�a�H�{�����ݹ�U�8a!i�u�d�7%�����Lsla��v����0�����o�猬p�7��;ܜ������H�*&��L�3��x�h�ޯ����|H�8�;1|�� G@&�b[�=����}�5�1q>..����&�Hc[5!��AO���c7L�Y�N�hTЋ�RM����V��yo�N�����}�0V���7}W�)���rj5B��/]-@����+J�r���sW<����60S$�G3ed&/��c*���QD����3N�w��?�i/�dd^��mʄ*�P� w�L�23�?ޝbC;��?L���6���g��	��t�$����+dhAS�ۀw\ll�i�p3 )�c��p�`�c|_P�ʢU�!->��ǖ�(��Sub�eǑ"_&��0s�"pב���t����C
|������ZЪ�ହnݍ1c��]O�r���Y��hy%��p��g�B��ðs��*�K���������E�|
l*>[�xu�*�	�z T��MhT�2��u�;���N��}���
��x���cZd`h����h��n�ͥ�^L!��y�#C}E�Q*���$�jE���ON��z�R)��G>��hI�S�qNۍ��1�=�J����;:�O�*��l��������_����*p��.8�]K7ɮ����R7�p�[H�^��d��Y@ms鍻�?9�K��ϱ;{�٧����7�C=�ey♾�F��/^��<��4I\U8&L���$$h�k�����!�]\\��r��|G�g����
���f��);ɳ�VS%��.�wI�:����N˵��,F\`f��]vqY�0���:����uؐU��A���3n��l�~$>oZh|��=V��%������ĮR��5|R��oK�(�m�+;;a s: }ј�����.EXxx���$"���9_/ZX��omѽ|�����0�uvv�������|J�20(�[�e'�Q���赆��(��cu�٧��-�)Zb5N.ޯ�C�����z�}�ͅk�����9̠L�㴈?3��5iϮ�&�$J���zQ��f�K�-{{�`C�GsQ37ׯ�b®lp&B�7�lkm�}�����R2�r��I�vtj���j��u��ŝ��gW��/�_UU6"��h��vS|_�HH�a�{tg�=�D:ڃہ��A$��k\�5�J�8��zT����fR�}u=Aӓ�����F����q�w���.+Kf�-�kj�/}��E(q~�qM����۾Fz��N�r�giN��g)&�{�w~F�"rr,#��,�\���푞
Z2�J-�zC/��<y���[TV��}�vK"G��T�<<U�<v��<~��8[YM]�U�c��՛��0��V�����6��ӏ�q��}y�i���6W�;��k�Ə�b�̯��x ~��I�X]]w������Y0�g��ѓh'�, ���v��r�&���MA��vc}�p�B���}�)yq�Y��"�Ă�<����yu��V��1ǵ����vy�M����A�Crx�t���pD��f��M��s�����0��<�a�6E�4v߿]]1�K�kݚ���۲��~��_��B+���ey���,���K�[���[qY�Ϫ��=ǉ�	�IG�����������9���qg�����o�&NZ�/X�h��*;8��_� �n��om�6'�}���R��Oj�&t"s�vq�S��c������
<����>y˲�0�d7l�>o]a��cz.�g9	��t���ݯs�y��L�}����%��\aW�~��6�|)((�6�^���厶��5:mvzǜ�y������	܎�y�����r�̼>C�Sg�����	������@5	r�T�����������4(�Ê�Z>;����M���A�'�"MZ�\\\$����٘�O&9_�P�
�
L�w��'ܸ+?��Hh<����,����S����<`1�gM�܆�2�\�[�|{�͹%����e=�,�|f�C!8̑n��� �������Մ����p��Ή�9#Sc�K\j�E�^_�D�&��-����>\60���V��3{YY�#.����]�/Y}SJ7VŁ��c�~�X^#�ya�m��W�2���J*��0F�/�h�C�Q=�±;��q��!��s����23Ԁ��ݟm���(.���F���W{�[���]p=[g;�*���qnvb��}�����5� �q�+cRSj5���&�*~g���+V����ݑ�x��(h�ܯ���m�@��l�"�P�$�z��BA�.���:����G�1�p#������YG�4�M̑�k{Z�uʏ��Ì��G�o�N�Ϗm#��k�}:���t�����fާ.��qdy�sݢ�����\���ԙ�!�;�ֵ��� �NM���G�l����l�pT��է�y��B�2�ܳ/�l��p�?V"O�)�ꅈ)D�]挎2��'��~b�2�O*�O����o�p��	��V�@�ſk��s�ju݈S�)y:էC�D�K��T9�J�����_��&DP�We+�����e����U�(� 뀏��5��@�B
�9%��5�\�>}�Bd��T.0�]���_V@�"Z�d�w`�߾0�G~�З���:{"�߿�|1c�7����!A��$e���W>q����9i���I��N >k��K�N�ɜ��-�������7in�^��1�{�<�����a�&��j.U��um��0=/(}�9=�(���B׺6͍,��F���ʚS����~�*�ߝ������a��/0����4"�B�j9຃�??���N�k�1��<�|X���~���T��x\���l�0G��f�o�'Ჰw��b<%K?_�#��]BY����~��|q)���&#��!�����j�g��m?����0`j�g�y�x��`�f\�OM�����ŏ�bD���{�)!�ǆ�~�kma,l6�O!�@�,�t��a�3W�Zr~S��4�@VD�c[GN+J��_���;�5��%��Ƴ}�l�/]��(�>`���_�3/�u���z��ƪȕ۹�n�	�ﰑRWA��;!�k�_
���|F��3.��,��/e~(M8��;���V��
׸'���qK�r3�Ognr{F�C�Z��`QX؛�{=���E���bflԄA��0��i5cQ��څ��K�A���^��\������UUUd���#WX�o#�<�o�J��;�)0�1��+���
����W�����*zn$.dRH��
	͚���AW�֘O(������c)������W34��=~b��2������c71����>}��oN nmő�D��篋�`��Ez"bVn0�����7�=�4�^RҷOΒP���)������'�����c�q\�QcAH���d��h�K�n4.
���v����_V�C�7Ly�}����U'��M�?2J×j�Ƕ(}���r��Y��L�X
�ߣ���}ꨴ#:+$�Fw�G�;�	�
l��ǯ���
~}3!���l3��HO�D�њGX7��;��յ��� <��#��XY#62�����D_��E�J��k�(�����J��(��f:�z�:�Cn�,;+6z�Q�i�<�.��?��Eo�Y �4ےd"�~�D�o�ŷh�?�lТBX������m�W�:m����z�^�n����d��.�^RYjU,�SXfa4�=�x�í!�Ĉ O�<~r���F��Z�a�B�*��ߜ_�ѿ��-��/�lh�9�.�(+޽�ɔ��}����#m�2R�~"r��m������|a�ຒ]�7=�0Q�C6C�SOy�Az��/x$�·[~	�����,�����]�כ�2K���m(CIS^�+��Sۑ��C���ZP��K�����T�e�!'�ސL�#7X~`w��q��:�X�y�{I�2&M�v&N�˛�,��ʄ���kp�"O^���D�Q�����m�U񼹩o��8���8�_{�T]KrG�T>����4%F�ոϙ�D���U/k|[D�u��(J�*�����:�l�|h���00h~xr��"*M�ʟwqqx��쭍��������E(K�|(j#JER�?z��m��\7T����"�<�a�jm�j�;�S�J5�����y%�^`S1�����������������,7
,~�J���A�>��%�5������c�y&�` ��Z�g�'Ɠh���	�ތ�V���p�`��+`oD�����܃d�}��"����8Z��D��P}{����xB��Q��7�N�g��[ňU޸�3a+`K�`q^.��V�?K��j��{6�U�t����kAJ\@ mZ���/=���1o.�.uA���
������Ba7>��Vmf-)O�+�X��,�����'Hᤚ�b�9[�ȟ?A�2���QfnE�_*�o�q�x)S��F'�cey�ܘ�E�	���ތg8Y�A��Jw((q��<R3=BώE�櫾�>���Ϛ@��%F��w��]�땄QGV��%;--�䥔�G�O4��*UBtp��S�ԧ�Q�g�c���>7ܗb<g��ɍ�����Ƃ���ք�0q!��т��&%���|	�:�q�/�ehXX{���8��$����n���~�\��fթ.j��=�=/$3���-�B��<�lt�'M�����Vf�7�-M_���&���[����;!����u3o���m��_7�
v"�7��aJ�ڡ
�CY�?u���J���x��98z"H_*�HX����Xt���Ta�f����(Xh!}�?����c���O�<��D�z���&rk��j6v�Z�L���;�֫�.O��c��(˧)O�P��Pv-`�j�Q��ݵ�<�e������h>�8���#�,�}ð4|�3Ym��?b�:�gАl�e�Ʀ��R!�Y��J������� S��M��v;;������!2�K6�-��4������/�n[;&�{�' ��VCCc��rQBRq`�����B��!�1�T#��𑜉��U�γ�3��C���k�����g���^���GXc��`�a0��8�:o��ۑ�#f����E������Dl��η���]��u�ip�0��-~9���@��~v�����<�A�'����@]]�E������LZ$�
 �B�|���CC؏�K�d�>lW4��6ţ�KL�-����<"[|��߇�����o�K��PU~���������O.��?�A�v��N6������99r�=���Zux����`���R�q������4��ԏ��gjj��k=t����A2���i�rL��U (/�ġ�8k
����%���Qˈa�����+7���;gg����@�`��5�p�ݙ
�/��+��ԟ�fg�����*�A�q>��/� 3�|��Q4Y��ύ�֨V ����@��S]V�4��
 ����o���ټ��{�O������9DE�te�o#�D���������cc�2��;��}O���������������������/����:����P���q��8�"����K��|,��f���~�'Ic4���#Sԯj9��ߥqo� �\�g��k�F7�7o�(�B� Sr2�cn�ޅ$�g"@M[���������n0��:$""~6��=Z��}��h�����{�	>8JO�]*A xv�(=�p���~hL���#"#?���Z�V�.���ā�ļ�V�7I�{��f��q��(p�/�����0��`�9�����+{��&�Ș܇�-*
!���G�L���ͷ�8�A��^�����f|�R\~�~g�俿P�y(��W��U� ����%뛛�dJxI$�R��g�Y�dX�bZZ�ݑ�������������<=����������EZ�a+}��]�R e����iSԡ�@�Qo 򜳳3��21�f)z���p����$��H"6���!���b��T���|��N����"!]���Mv�M�����AEx���.i��킚ņ탼�fS��3ʷ�LL�e�����O����G�k%��?Wcg��7U���&++�*��mP���%	&�����σ�ͽ�z`Zx:�+X���.<�z��ن�w��2Ʒ
C	����E�^B͚��i*�����Sx�1�s����h��|�Qj�e��)1��H�L��8�"�Y���+{�.��1#�|U�R�Z&��p��n�u�w�j����^6`6Z�1mnӁ���2����H��)@�f@�l��f��'�Jԗ,f���ڤ��냟��P�Έs��7_G����c9��V�Q�K�������J�*�J�$���О�+�G��efF�z��aܥ���$�9��:���U՘�����E��6=n�o+���M��,���+M_1��آ��/�5@y.�۷eh�n!���%s�>�;P+h��ٹj��-��Y�V�=""����2:86/>>>#+K|���?ө]���Z��"6쮝y�^����7�\6OmK��������Z�D��aI-hN�ߎ/������ө�F9P����K�,k��>-y�xP��,/�����G���L�h��hgHZ�7�±�Ӑ}��=5�u?D�G����3�9m-r�=3��C��-ǋ�qT{�W@#��f|�8��� �}�zL��D�:t��a�?��f�cb��������O�Xw�JŞ[pu/[^��=#-FBcҿ��iֳ�p�٦�hT�ت������P�=hoG�V��꧜0�cpHIC�w�� �b�6"��� ��I�L��e��)ڥxe�/��������Z�r1GwHiBr=cf���,�NT�g �����V�~xx8��J]B	["vvv��ё��߿�J@@6�I_G'|k(�N@�����8Ƙ���:��"�w���R܋�Ey�U#�q���Q��B��Q����-�!�`'���M+E�����TR��*�'96�Ʋ��SN��7ym�/�����rW��
�&�r����!-j{qI1!>`��ʡ}=�TT�9�@C�K-�{r�>�I�3�i�a�F���k��;��Wx�_o9�N:J8y�ӌ�rX�7��K���-���Î��^��Fb�������˹r�~u��Bn]H��K��W�+�ӃueY�[���ٔD���0e_�{f93�L�u2I폭O�Xrw �fdP�=�r��%�,�͑��Jn!���TSSÛSטZ�W�$��d��:�ae�2���69K��4�U�f��%����z�#����c%�>�h��f��������z�|����1�e#V�Fݒ���P'���-:��5�ؚ>��d<�^��D��]�gO����,P4��.���*��Cx�eS�,��{�`:{i��r��|��9˖��$gc���@�U߰!�g�����Q���_�+yy�$��j�b!"�:�~4^s�c۪�z��Ք��s8a��k[�+W���[?S+��9����̙l��z^9����� ��{"�]���^�F�x�r����ܻ
&z��͸�P��gñ���W��&o�M�������8W[�B������C����ƻ��D�TT��=<tI#��!R҈4Cw������* (����0� ���C�������Y��p��{�y�����9��q	%��&&���{�t�g,�N�ỰjmF�kL�T����S�5������a	w�Aå�UWW���;����r�_J�!����s���vx�h���1m����7���c_�q�
�͛3��/_�MOGVTl������=��UK���T�d����MХ˩02�.���E`5SqyI\��X����[�G�����z9?�l(�Z;�uL%X�rB���fc�?T��9�<�}���Ltz=gZ�b�����PU�x'�$�����PC��zb�V�)S�"�Fe|6�!~1%L���"+T���I�qis�<����^��Y�S���s���?�!z��l-�5�Y�y��~���<�}	���x�ω�O��=So�T.	-BAA����[K�O.&�XYZ"JJJ�I-,�oa���@dd�sӖ�a�}$\��]3D�8����󍴴�ˍ���ť�ɪs�}�2�m���u�&CFC�ܟ,R �@{��`V����l�M`�m)���������7��߿w�!� CVS���Ѱ��2�L�ǀV�� $ ��w�
U�xB���Q��Q�[���6P;Is�X_�W�]�wg+U��}U+��O	ܜ-:S{Lv_�&�̰�Ӧ;�W&Ɨb�ˆ����k�{LW�U2Z�d�H~�N��l���`��3�bF�J��M�k�ۻ��ł�Ym)Ş7[W��;�uj��l���|���ĝ";���-��0�}����~����iG|�*ˁxr-���x��7�Ar�nyXBB ��H��d8��Z�mk����k
z|Sa�
7�'�����̓���{A-�	�t�=�����{�>�gh3Cșxy��
��n����SOnMALL���J/��U�n��W�B!�o;����C$�n��[fq����Q����r3�֛VؾdW�ן��Ĵ�1u���&�-�uh@D�W�C�}`��QϪ���G�t�g�%Ŀ�f�^����ID�zyx��)�:v"nX�3+nek.��{���zd�h&ɫ]voβ���nY�]�[���L	2�K/��a�����͚� ������@j}/���kѰ�9�`�h�0�����,{��I�]���q��p;_EEExD��R_\^~���9�'L�����eac�fcc#,*�#
ٛ�f8::J�����~�jRK��F���{!+�#L�ä��N��l���<t��l���G�Z44���o��J��Ĵ�U�e�蝿���t��$侧|���^l��疵Rۉ^ߺ��e�Ӑ;��V� ܨ0=� �ո�ױ�U]��gSc��}i9�!3�4*�kdC�~��f���fmF(Ὰ�7=ֵ��$�����>0����Y����;dDJQ�����-dǕb>��ܦ&�Հ���_��`��اOx ��G�5 �l�G;�Bv.8�����S�LA�4�S�Q�KRy�*��cG���og�.�!#ҥ�,��PVn�q<��!�ђ�0�t_�/���k�/Ā}����Xv��Ė�O'�j����:g�!
�����tqA�$�r�D_��533+�Q���F��u!02�6�lJQ�L���N�p����쾋s 1�蕬��'��q>��^Lf���>o��c��&��ݴJ}hx�Lާ�rk�R㦨n ��ԥ��	�p����x9f�稃A�gyݑ���ux��\ݘ6�ϊ�JA���
�z��@���&w��nB9��ʺ�ą��<�����ǹi\*�`x:Y���?��usmw�d	#�_
a����p4|"���G)��v��j�j}�W����\t��z:QM��zFe���X�J4�D�d�=���%�����J}^lo;%fX�Ş�ZD���E�h��YV��H�$�RW�|�V�ud�Sś[��� Ȗ��I�y�á�M���|j{A/�@��W�ߗ �F))�/`���~>J����-�DXZ����je�AƳ��0�.���s��{��]l�����N�13�5:��q�;8����0��%`5 I�B�+�D�o|R
�ʳ�7e¢���g��ߪ���:>9#y��
	)(����fT�_��!�H[��Ӛ/�gQc�C��{�Rj�Fآ���`h]�6���e�
j�ZϧSb%��D�/8%������[�|9���y]DBA(�M�{{h:�zӀf�-�����O5�q����G�C*�l	eee�>�^Eo_�索ۗ���SS���8��h���FFFGs�0���r��)h�jD��$ )��f��}''�D��'�f���@�&!�p��Źx�uu��Ա@���r�-}�o�+Ģ%��Hy�k�����Vx�X#�5�b�O��
�;�׻�U�u�(��6��~`n.s�=���)�A�>6r=�c��VP��H�5����н�{~�E�I�gGlM�B6	�d~�Z��AN������ o�DDG3��Q��]33�Yo<�22(2���%���`�̕�fUSi)������Qy''nM-�ϙ��pq{W�����&_a����`���.->|��)ӥ���<T����n��7���W���4��l��f1���l]�@u���)�Hˑ�g��}_
U�����qU��'��e�ND�Km"I��]�H$�S<��DCE��[�ph\z�i3ܠ�Z��'_��f�=��㩘�c�2*�r��0%U@����/Ǐ��4>��O @O�DRj�D�����.����3��].�������ʰ{_*d��Q�6�O�p;E?:�C�y��!�|�o����ҫ4M����P⠽{���=&�'go
����a�F����'??��xA��������Yyx�a���#���;�uv��Y��Q��<��<�,,h�_9�������W{�љ�ޮl>�3i�{>2҉Yjwf_��Yk0�_X�E�S���F�b7�?���P�֓���š�S�Dl��k�Wu������ާ`��<\��PJ\�9(��L���-�I���l��+w�]4wH��ـ�2���&4��MnB��D���l����;�#	��H�~R�gj/�g�t�};����J~�E��YI�o"۰{;���b�n��1A����/8�������(��|&}���Q<�u��H:�S���s��bX�MM���%�f����vcT�9�J�,,u���
�*0��C�9���s�3�z�h����0tc:�0.������N�?tuj�������M�����c�@��Aޡ��;y�+������L� y;u�W�}��i"�_uo|n���hT>&y˷�?�rk�+èxX�jѠ�6�Y����^��{��ebFH�y���j������nL �~'��V��
*\����X�ݖ|�Cxˢv�/�[��dv!H�PN��QL}p8u
�(��M��P��D<� Ǵ�eF���;V�J��O	8�{��~D^ϣ+Y��z7a�OA6MoUK5u�r�^0&}�k%��} �x[E��JwE�E�K� �����$�<F�\B��O�	d������b���_��(���\B��6�S��=v�O�oju�KE3W+���K:!�����%%'P'1Ȝ���� ��tsg�;�vH�#�'`kף��6J�g0I�xAq<��)��&	<4��i�����~�6m�c2m,����uȕ�\�5�E��I�\Z�\�b�Q�[Q��ҵ����q�=c ڬY;%�K�DT�ʻTmt^���A�7 ��ڶ���}h��g�5�ލGEE[]�]M�jR. ���ġz�z�9���!Iс�GQV�2���qqE�N��%G���c���mk>|�o����̢�Q�z6�^8ly�
��E-��}��?�8���ћ8V��	�-&qV,�Idޤ���G����Ҙ�v-����M��$`��Z�Tk\:z���q����a��HB��'�����U�,�X��j�Uu�ڿ+�3/�lg���2i%�^�e�8�n	��¹�@Q�Z��Iz-}6j�	:*�f.��
��H����r��Un��<=�Xu�S�4h��4���T�K�T�W���K��:4�'�R&��֛9T���#Fp=�Wz+�E��V���@c��[$�O��ԠT�R���=�Z/�Nr�w����9������σ�I�7t+�cp֐�>R4|\�lzKO���C��~�����������-2��������Z���{�.^{<�k�$�~��g�L���{�?3��6I4]�Վ��5�w����?\F�)Р{L]9���P��=ߌ��wl�:y��y^��l�l �y^�X�(���p��z�O�������q1G4*��<J���b��E�W���H�����\+
�5�xNm^(��{�GZ���s��}�n�ڛ��_@Xv�#N����0��ؗE�������VmL�߮E?!��rJ\��D�:MV�SX�2$�ä�����ۙ,�nSǹ�$�sJȑ���ctT���h05���+��p8S~$�"��s�h���L9�v�ˇ�����d2J*
4����$#��C�E�DK1B��J���[�έ">qT|�Zv�����|뿫)��5���d�Tޚ=AG7q~0Q\`_RKu�B'�ԫM�wM=�-�u��/�I����EOV���<�`�gg�*T|Ϫ�������;���F�M
���l���nɮ�P@�H�1,���r�l���p?���Dё&�˝����OVbw[�>��E�Gw)j�aٜ���E9��aU��U��ݠ�Yy��MT���h���{���i-��ir�D���/�]IT�̿�;�+����Ef�����5ݷ�ə�@���_�P5�
���ǿ000�,9�n�v��� E5Wm��p�H)�j���H�k��I�Gg�@��������N$>���$N�H���/A�q��@0z��������	�v@�+-\\��_Mf�y�{N�4�����=���]W���ލ��B�����t>$�� L��S���� R.�Dῧ<8��O��X����ft�Q�����~9�w9�-�=0e��9���P���lu8��y���m��?g�M�% �(��Ti���pt�h��1O��2fEA�<���LB1�c�O�[�F�o��r�HC�z4_���w�e|b"}V"_�h�	�~��	B`WJ楘bN������}������4���Lɻ�ը��i�N?�� Gy��Y�A)\'�����4��D�^X���Ƣ8k!��
9θ{�ʹ'�.w^�����Mk����?��9W�]��8,���?m�<a2Z�4u޺=f������o�)�~ <�����Y�N������:y:�L���;���q�� �u�bc����ȏ����4Ϸ64449�΋�f�9Ӽ/�uo\a�p�T��8���΋��8p��.{���;��V�!4���D�}w�|���p"�ވE��ĭ|�i��e�u �{*2��=��0H����e�j@��S�>s �6'K��F؅6�%�5A>��;�)كL~��:�b}]y�g- nS]�b��j����Pà����2ݥ(����d|v6���n��jX��K�˲���z�$���&Q���Bw�7>�1d����b㽿���������� &��h�r!+q��teP���Z�&�q��t�i�WL,>@w�f]X�O�����c�`(���I'��4�_��1�,���x����-�'x�_����JYO+p;r ���؄.E�Q� ���J�2�F4�f��A;��M;��K���40t���w��Z���?���;.<1+�o�q������Ne;���&�݄���W��k���SAn�I	Ҳpd����*DC6�����+0�઒Ř��&�a�����Y�`q��W@�����`���Ï�|��&���g���T��P'Y��@�=�~*�!C�b�r��^+���"���q��@*�}��e�����^̭�Jd������Ir��n��YN����{g	�����/Ͼ����gk<S6�T�셩�3��J=ǉ�G�iv�n8�Q�@g��Y(?�^XXh��v�X����Ǩ�8��=��Ҳ��y
B�I8jE��ׁS��.���Z�����U���)��e�2���^'K"��p3E�;E@�{�K����`�	5\&�����Yq����L��?h�h+�2���fL`�S��^H�C81Q��w4����x��PBs�cJe�6����`T��a������8�_;��8v��z�@���%�2���w���7Z(`W<@Q�;X��3����"�J }���&���6��7��#��*Pִ]Z���b��>W�k�*���`��;��o�y��b�whŦ��V��S.I٬I�ʓ��� $h����b��R����X<�9-K���4�<�7�����di�9�s0N/�,m0ueDDD��o����a�R�p�"��Ңu!U�Шi�h��� �>NU���^~�C�,*ﳧ����j(L��K��c���~SO�����i $����>�� ߖT��2��@w��<�T����(�� /��i=�VP��ޞ�y�"����Ͽ �&5��0b\T#3qſG��boV��¾xIW�{4�����:V} k��V>�H���w߱�=�i �AWdb�wa�<p��Kz{�Ҵ��t������V	l��!�!����sL%��p[!%0!��$L���W��/j��k�J^�Z���UL2G˱y3tx�z�v~�a�2����E�$��i/�3��#ꙺP�0L��*|hC���URB�/r=���ƀ�-�]X`sj������m�0�@�&y��	��������o�ʯ�e��5�/�H���{қz" �a�� %h� -��:��Cj�ΟgIJ����L�߮�
E��"�\n͖o�n��W"�*łg�cz��9��O�0�ʏ{�:�Ʈ��r��e�@�y��T�%� Mu��:,V4�CVE��_�Q�	W�~���!����E	���O�%R2缢@��*M������B`���[��1<(e�hD�������y����j�}=�yl6���|J<%�- }�TA'fȍ��a!|B�(�+��A7#�^�]�5����ހ�9��K� �v(�kBc[Ի*�_�F��&N�u�����q�w��A/ ?��������2�`i@� ����`^�c������L�O�n�x,��f�V�Bb�	H��?�w��O��#�+�Tp�8%��_U ��`�V�a�B��[�f�D�X���PưD�Ɨ�!�SgF�N��:M���!-�H�%Ox1d+��ׅW�s�=�z���EE��HX�顪���:�޺������k���.��f���G�B�ĩvA�>�o.|o�µ_Qy��dK}�_4��k U_@ОʠR%㵳豣͌
�TPv��|%<mp�w�*�WHGq��Tn��D��j���b��8���ߔ�XA�����X�yږ�kx,h�}n}��dX�ې��f�<��?Ru�};��Aw�[zq�s�䡶d�Y��)�Έj��� �����败+ʀv�N�pAHO�����'�ɚCd�-�V�0����~��?W�8d����Gd������-��Ά�]�]�d��K�b6���x�;��>2��Q����X����di��Ux��zK1F�%"�a�6���!3�";��`��2RH���!yB"��6��2�]j����Zެg{��1j�d�:��J�5	�g��)�Vu����&2�rw[\~�����u����Ah�v�j�z8��G�g{���J�q��	�B�&�����D.Q/��/RV|P�^*��;�^"��	�Y\�j"��]��x��9j�D�c�2F�	�WY��[���k�!Z�5kL�	P�#�<����<�� #���"M�"wAaB�����UVT�b�e9kg�	�E�K�����~O޸4�w2�����#13��+[y� ,&|�.�a���������+��	W�
+*�F���N��(LR�����\������0��,�dGH�\��
!��#Z*W�%o{��u)]V�Y8�b��@	���e��.���a�n�+B+ ������M9Qo�F��&5ayoP�����h�9�F=��%���젧�����Z� J\�+�l��b�w���;��']z/�n`�Si����F�o�;~�P`*0�z��T�F������@ aoߪ��hR��b�����{g�64�A�O9�Q䊞����~z�ݲ��ȃh�a��-u3׉�탛#h`�QF�H�$��V�(�A�I~(�y}e �	��e/������G'�1�i�w$�Aޙ`��M'�phI�|�[:z{%;[l>���|_n�$q�A	(2]f�	�	(�de��.�k���#UK7�*�O�"b��J�JdN�E|�,fog�T9gt�#��QV�0�����J	c�ij�]g����׮��'� �e�H$�R%8X���r����&N(���帐΂x�3/���֞$q��S���� �9�t΅�9��b�e���0�;ի��v�&��CޥO��%��Eϼ�g]n{����G�s�k����U�e_���'b�������́�*���Y٩c`��yI��ߡ �}ˋ�A������u��{�w��QT�:R�P�
#ټ�S�Jm��L�=f������&�H)~�Z����C�̉'e� �	|?��\��H)d_�����"i�i\��?����K}��!��t��;�'��Z�Kt��1BLzq� xl'\X]�T�.0/�B���8=��h��oaZ?&��O��������aL�|���{������jO�+n�Y�j3"����$qO�ջq���a��1)�ƕ ��?�
���s�x�V �{om�ʴ2�u���0ȗ�	���Z�Z��9�&9�j�m%�MAWD_�_�x~��eu ��雹	dWD�����5Ư2��U��A�o� �a�*�Y9�l��堐�e�!o*N#�M2���-k
�����)���A�7�%�`�ƥ0�����O
;l��ЛӁ��+&�����0Y����g\F2uu |w;��o��S~�8�#z�/3:�\nB���h�%5|x|��:����1�ͺ��o��/zr!����6�tZP��o%�]my�xHX�Q1�.��]ڨAD5���[L�_�cYB7����q���"
b��c�9���f���J����f�{����@�&J�!6��	EN�(��"��d3�KU0��0C�O����@u�5�|[+	�m��%?uy��4,d-�����굻�E�I�̀d�]���sv��Cc~'�r��d�;�Se�m�V�2����+�߹릣������(*�s��o�qѢ�f�]��z���O��s��	�/<��
�f7�9��[�:��nT-���;�ǰ'���v]C�?��gV����Q����RO�Ώ�50��B|��$,Α��}H���eu1.�"���FJ���K>3���B�.fr�o�=�*���j��S��	\�G�檳f�[Q����&?�9�o���nv�ߣ�f�\Y��[��w<v3,��ba�:)��90{���H�����"�r�:Dl�1�(4�(:b��������q/aӖ���t�`z��RG�:�]p����4/%�+�U 1� 4�O��0>���H{��M�qs�֬p^���c)VFנ�%#�9�����1�䴧]�v]����L������9ͦ9�������9@�*lo�M�ӄ������Ɗej�`6�O&.�E��3^R�n��0�� u�Ȗ��C��bo���P��m�u��sǧO���K����.m�U>ɋ:�ϼtĩ�k��˯�������Fo��]��P �)�uw"Wp���i�H{�󰕬&�դĶ䳙@JM�vv6�M�8\~8�O�c��\<eX�6��s9�lkKiI�ɾ��Ԏ�y�wJ�^���9�69.���o(f�Z��-O9x�\����]�##���}?=Ɓ���:���L����rfm�x�7` �ʔ����-7|�M*0�{�yR,˔�g��p�-�R̳�=���}^zJE��M=p(XY��(l'��Q�c��F�B�1*���֘��kN;JVU0��Y���kwB�7���-F�3��	z�k�i��U����(��B>�\�Ǉ� b�"o��c�����7��eVd�C��`��p\�9X�ݮ����K�&l1�Y�U'�b;�L���z<�3�t5����iᠢJ� �r�_^"o5��`w���Y��ܬ9t�C���i�����<��aci�����9ϑ�R`<�B��A���wbWco�Mva��wJ>�	]��N�떷#�͚iM�� �$�eZ�*�o���}�W�ۜ~���7Z,<X��Ȕ����`�I���N����$q�B�mbN��ÒI� ���_���5�"1.�gMQب��T%:�֋�Z3,'�UAl���f��|�\b������<5�|�Jw�j/y1����#[bxk�(��=�$� m3��A�D�����Up�3�ݛ���t0�8JeT�^8����GK$;0�s���a�G��,���N�����415"�uM;!(4bR�I2�6_cS�M���f�?�E�^�H����n��y�&I�]g�&'կ@���/h�afD�*rӝ9%k���C�ψN�{��nh�y��ui2��T��s���C*B'�ۙmjy�z�1ǸW�7�-���r��T�z]q��	'y$?�w�}�r�t��x�b����q�}cҔ5C�0>�Y�HjeQ�G�g��&UM�?!z���ԧ܊�`o��޸���l�T��F�Ee8w�={�6n�����&�9�9S'���w)�������&,�{���{��g��C&�(to�Y�:���._��o�,P`�GƂ��N���82�dm����sl���*9:B��|mC���ΒWu�bb�/�K�-,�X���p�ֈ��m��;#pls4Y��k����>��w���ӟ��z�Z<�\7�ĠG���2T��lk�[��/��(O�����PS�yt��B���?���d0�M1�0w���g�4���h��Na��ħH���b�#��R�K��? ɒ����1�މ�0��BP����$.Mܑ�t�%;P ��`ثj�R�b��)�����q<��-�n���^Jv>��<ϒ��ǩ<:�,�N�l�$-�;��y~���vx�!�1��1�q�.ûT���}�O dڊ�QQ�	�8=�{�읇�lwi�kTc2�/��j0��%���ݱ;���bp�h� ��Qx2i�&���1u=��Ty͖FY�"z��/r�{���~�`D�F���I���N�\�A0z_�N1'���p��$AH�>l�c#�7a���4�)�G�{H�拋˱U3�mg/ꃹ�7�]�e<�Q�Y�D�W�#��8����d0L�m/[���V9}�y:<5[����+s��e5�C�}�[��}�_��U�FҢԀP��A<��4)s���������,�`�̫W ���G�	�fqM���%.��0%�\|-r�A�1`1���W�%���I�M��兺Sd-��#z:�%&��c�Gl������>���������#n��K�;�����xg��ɣ��-;��@��ı"v�
���^*���e�����pVT�D�,Y���E����CLa��y�[Ňi�^��G߇���*�-M�V��}o�߲E�K� �!ů�6�_\��-~�拳fq�0�uUK�ԋ�'Ǖ.k�Y�k�p�n�'&x��L���S����*ns�	7%�ؾ��.˂���D]-��%��A7b�u��=Brt�Xn k%Z���zО�ΟF�~�������hg����;�ASc����7���]�#�&ɇ����c��x�BJ�a��׍������'1���,��i��HF���BM�f�3��T�����p^��.�L=T�I0I_�����,��'��B�y��fa��jLh�4ˣӂP� ���N��'�	��[��
cs<��h�%z.kd���sM��a*db�.C|�����(��j>����%�^�,���
���Tt{	V*mkse���<����H�b��Ao�n����뛱f�7�:�u�g)��$��
���
�C<��ꃶ��T*������ �\ ��8��������s�s�����k?]�>u�AWT$ʩE�XJrH�i$�?��,E$,��n÷���ҧ{-*2��l\A�b��#s�^�݇q�e�ɇ�����0~=��b���O#BYُ2�O�䖣@j���	7�/�A4�R@��6�H��|M����6��^�ͪBd��O�z��F>��%��)L[l
Ή�e":L�4�6a������@V���1��c��xj���fRV�4��ߠ�=-�Tk;��>��-pYY"
��[����N4D��It� )s���洒�T�:첍�J��*S�	��}���H.E_N�n���	_N��iɛ�͐�"���,T��w>�i���Ǿ7�rn˖릠��;yp(޵[Wo5~��j�2G�����:/�)��@�+���.��t���I�J4#*+.暇�������Y�w���k��%�J{m�_̎�l�A`���TJD"s�5���w�$�$����������9�u�R� G���P?MSV�2�����@1y^�O�^�m�#%jb��(U�0��Zӽ��@ [�f��'Vd��U�K�b(i�Ҭ�i����e�h���0k�~�;'���O�@��C�]��M*�%�.�&!,��"����Y!�(�����3���T�1�ƞl���T<?�l��v�K&]\�fLK+3��Z>�Eξ�1��bhqK;�%�G�w��K{��r�ʗ�APEg���hC(��B�@�c�*���Q)�`�G'[����q�(0R��MV����XD�Q���|�C��~G�5����Q,#a��å�x�Pd-�6k��!�.��H�]����(%�Ñ���:��v�s����h�x� d95�NM���\!b.�|a��G�uҁ'���%'��U��`�f5Oe�N�}������6ᗓ����k�K��>�����6������� [[!���٢�;�G+_0��&� ���1=z�`�gZ�Vbn�ӕ�Ԡ�o�=sb8[1�/�
�N2�������Ue�q+sB�d���V����u���W�S��}�;cG{#k	`��T<�߆upj�턞�R�#S:P�H�/�?H��n~�[h)ġ��k��4`Wt��{G�q���|�^���稄�5��ѷk�LO�)��"0����.&w�^5!�w�\�	�e͍��T� X1Lr�D�cӈ�Gb_���oߎ��������밋�|C��#�>��;��եE_t�MU�JŲ�%3d�H���Y7��d��%�$_썈�����|����)�bo�h(���;�
������NK���- g�юX�dŶ��Jy��w��f.nn�s��tN}������@�wv����7� �l]��ژ]{:��
uz�\J>�>wa��G���-=_.�)^�opZo�P�#��Sv�F�!�o.0������&f7��@���mą�������k���Κ%� �DeǄQ���S�CX�̢��K�I���O�H��(�ޡ��� %���x����q���|i��	 � ,a:��H�{:������0}yQ�yZ�	�-�]����7V���mF��Yb�?�q:��_��M��:a�-r��M�?���q5�%�'�b��pѹ�
~^nRwwwU�6�z8�m�㱳�Q����y���BK�Y�eD0X�-�6?��u��a�"v!��]�4cز`o�V1�f�����T����&Xv,�
��~�*�.SJ�[V| ������\��>�SX;��kRFq��>�� �K���+Nk`ф��m&�lߗ`�F�X��Q���d�7.�/'�	�L�7��*��q$f�l�>�G�%KI�}kL8�h�y>�|l���~�����py����n{�`M!��5����cj�&{ߑ$z�F���t��ė{�v�n:��C}�[^���}��&+�63Lv� ׄРl�H ���Z"�ۅymԬ��K~��tw�ed&anе�G�;>��ǰ٨I)ŷ�o���/����">-�~_\���J��eYh�5"й<�ԩΥ�
)I�|Ez�қ�X���K>�D�"ʥ���}-�����;��g	Yk�`
��xA1Th�~�W9�r����{{e�&���A��bmYB�# �"����z�@E1�5��ap��r��9k��+�@�P�����IW�N�ث;B~�T&s�i���>nZ�n`�L9}����i|����(Rҭ��A�)�FN"Z�1=?1ZA�q�xF!���K�(��GDEe�#j?���H���5�GCl@(r��Y� �I����r��ݕ����v�ce�"��y�	3�r�ah�Q����R(ؠ ��o�6��&9��w����u蝜fD�|��<7%0Siֹv���6�-��ff��H%zV|_�mt��0[�q���9eBX��h*�h�0�r̘KI��BT�����Xe����{���4�2*|����RyU�/-���.k���`�.#
�-��f�;A���O9��z�5�6�'�!l/��f�^)G�'�F������`��cu'IF��j21�u^[�.��,��	��'�RR|��t�Nu�z�y��`K�%�p�7�'x-+��8���9㍮-�OJIs-P+���wm�h�H���4ǠMq����t���e���J^��5������ud���e��n��/��]�'R�J�DI�E<>XP/(v}t��p�~\�?�o�c�� ߜ�Z�X��)�)ɧ��ӗ��D�c̥X|�jA�o�ܔz�rPHq�ݶ�~-ύ_�/�C��Jt�'9���T1�=[�ѐ�.ū��.b�AdF
�֛�пT%��o���&k��-vi�)vr�-:
�N�s	{ν?�d�>���>5������ {�Ė�_���Y�".����-�s�Ar�XϹ�XmA���Ҹt���)�ж�s^�s5 �|�o(|��k���M{���8�/�&�y]�py�ȥE��$�n����6ی�T$�o����w�%�U�a�L����DO����}��۽��	�1���Q��"�`zލ%���՜ӊ��	��Yܐx��?[�y���mKA߆�dL;�6#��
*�Pn���/s��`�S�m��_M����V��@�,z�V{.����r��u��p!~a�얕��hE��z�)��.���OxG�.g�C�/�b�����F�Q~��ڬD|������i� ���A����!�2j�k�	b�6D��3�7r�֫�j�Ք��R��t.�M&)�4�+����-R�#Ď�a�z��ӻ�{[��P�/�v�[!ç����,m��E������t���"����#��=�`��ۘ��=Q��盳�Bl9�-i	� Yr�%���$��y^f�������q��S��b��dy�	}����5����Gw���j7Q��T�O�.�����p��T�y�Bdc���u�"������̛OdnB�N@���싙
�EH��B��:,u	�`��iVc��ɾ�WϾ�����~ܷ#�7��&�� 6jSa`#�M	�
ˮ���^۾��TQ@:��ě��.�_�J�cN��ޓQ0�H�>����*e��˹m�i륇ia��Ħw��� �FM����H����|��G�)+�r7�>�Ү+�&��T�6���s�4��x��n�ױ�L$^O݌��ux��<����N<P3�����t܈/����� זO���5A(���uzƹU\�Dɚ�X��=�2"��~2}�6TV������[�	�ƌsb�k6W����-�M.(���R�j�wCt9��	J�*.�÷��}O�"�8�K_�ms0&Sr�^�n�@D�����W=h�U(��)�s�Ӈn~2�+Q�� ����}���� �ֽE���K68�T���1�_�����pJ�)���9�D��<~\\�V0��1���&+�w��Z��[���Ǜ͹j+ׁ��1S�?���=��ǽ�og̊�9ԡTU?���-�'���eM��x�F��=�{���sCJ���q �i�}�����Z���li��oY�D���1�a5Ǣg^g\IT}�C�Ջ�H�F������]���,���i����/��s�������k$���1�~pĝ�+ޝZ�^Ŭ�l@QKD�&7�N�x û��o��f{�SS4#���K_�ǳ�5��f��(�x�4�Z�"cm,:����F����"=�����Q����1^��7⧾�����pr����	��
�=�N����˂˸�k��ݱ��� nK�8�~��+�*vX�S�����5���E�*6�H���Қ���煔4*���Z�@\��'��Ƙ�i�����uVYś#:��e�)�&/>j�@䔂"�,UD�.��H]��c|�C-n���%*�tj�U�An��6SKչ����p�q���d\����4���B�u�C*&ߑ`������kv����8�- %*.�n���h�ʰ����S:DA��iiDZ��Z���A�i�s����%��g����u�}ufΙ�����|�~���e�^V�q�����K�gޗ�/KH#ǁU��K̋�%)�T�����zΪp�Sr�f�g+✲NX���;��f��#1���Y�dPBd>��Q�?���Y��Ql�Cu���ޮ$vl�Uj8A.����������h�P.��8����|2'l�{��Ƈ���m��Z�)=�l�$�`�°�q?[�5l��Ҹ�]��EW����j�̺D�̜Z�Eh��~d��&�]t.\���3Q�U��E/������l�|�=¿�����9�ո�Q���uT���t7+ƼW�/Z1�֑krh��??�`�����CYWc���t�g?_����7\���kЇlMf]l�G����9*�\�Рƌ�ǎ��C;R^9>_$���6G˼�=���Q�g���V �E 5�B���:�X�;�21jA}�$�B�J^�T� ~w-� ��%��s#�_?u�;���9NK�j@�(U� �}�4����x�"7�(,�T@ĭ$=��$��t�>nO�C^�m[�����R�SQae�t�dQ0m
|��(%#bh�>0W^��@�suYT(��6�	[3Cj׍Jx\��G��ãڤ�����D��a͝��2u~��vI�<B��6���0Ş�)�g��|�8y&�P��K���C$fΥ�ї��p�4��KC�����Ix ���h�80e���ЎP��z$�q	�%��)'7�������Z�������Ĳ���|� ��_�v�G��FSǿ�����K���%#y�*~�˵q���У���C*�ǂ�L<r�.��8K�c,�+O�gBZ0�O��gr7���9ə�h��I��=m0R�ٱ���v�Q�l
�<�-���U%yyy<HU�]yO�����|6rkE�y%0��L�/b2�E˫C��/^}6�K�2v�͐Wg����w���U��E�ڴ���*�:=(X�ډ�Q,ݐ�}�Y��>�r萦#ra��Tb�d0�d>��#}.�&j�᥀|�MF�,���� _N�CHH�
/fW�c�7	�߼������2�?x���@z��32���ƚӅ~FQ�|�+[1����ݲ�?����O���M}�V��c�e���#WQ��2{S�?
�h⦅ �<("ʷ�*�E#S�,^xXS�tUvc�M�q�|����@H}�����x���L�8��&����G�����IK���6�U�-��џ��u�4��V�����E�a�Z�-5�0��]����\�`{!{!�UC/y�u�����T����Ϥ�0m�>x)X�ԇu�	�b�
 �B�o��6Jx_�r�= ��5��ļ>�����)84�G�xGMr��@�G�Z��E�C�X��ԑ�Ԧ&�E)7kW)�Es��O_N&�ܧ �ՐY��M'W��x��EI+�%C��`D\T�w#|�S���V�l��_�7�%`\��h�h}g�-�DFC���Ʒ!-��D��Sy���ݺ��F��#7�ߩ9�\���AF���� ��h�5u���,m叚0Ym�v"��
'E��.c��[��G_dbF��e��b��9h�i��H�������l��M�gl합���#��}��D��������#h��W���5����+E�T��$��錺�?��֞O.W$��_�KJ2Yx?�դ��R��]��h9���Q�hm�}q��v�U檥����W��7vI�/8;���0�����]7߆S�%G�Ք@�)T�a��h!l�w�J[`�����7��@������W�cۨg���
�hX�|�>ײ��W�!3	�@C/]���PUF_:�KVS�	X١���Ax�R�~��yJ�HA����_�@��i�a�(�.�����<M=bi� �έ���m����@c��������ԡ`ܐ�f?���b����	6'�r'p+��l=�ڴ2Ѫ:����r�E����@�kk�ݺ׍f�'c錒��>�������I��m0�*��d*b� �U���O�=����m|���%��d�����I%n,[V��T��~h�5G>\f,~~[@�t"Ɉ�s��\e�����ᴤh�vUa	�]1& �"x'\S�Y�0�]��o�/�ޛlK�	��	���A�ehy���%�J���E	V�*RnŌ%I2�>%k�@+&�i�͚|���Z��ְ��F6t�G�U
ظ1�;�V���:�cn1�[�qm����f��W��t�,KC."��|�N�,����5����q�Ör��z`�?�ä�Y����[q���o�3��5�NB��9�1�y(�6�-09��8c�S�>����Ĩ��]@�X*��,�Jס.F��S�I�D�Dr�v��:+�}�_�(5\�K+��k���jM���O8�H;'45.�o���Z&��Y�f�F$�R��Op�[�--���$���N��s�<ˬ��1i=pџA��F0���wEG�1�v�{���Z�N����ٸlޱ�A�����(Z�_q�����q����Z�G��]��:t.����r��rׁ�����,���oF���������C~3��,�l��CA�80{�F~�05X|��9�Ϝd�:�Ŏ�5��9��Q����m���u��L9��-�(	wj�}e�-oq�~����H�;ra����?3(�-�ErDz����cs�`޺UU.������ӕ#��5��'�n�+�����μ��뭭>��O���;�[�/�t9Omuڞ��E"3O�^������R[iG��+���_w���?"�����,��Y Y�=��*Q��'�	c/�����0�/��{͟[�r1�Y[��{Lx� �#�� �l	M7��i��nB�w��~���8uM�g������B��8�8�Mm��o`��JU�.�R�d�՜�!3%l�_�|o��p{]��܄\.�4�=�@D-X�p���w��b�ee����""���p�@���(D�����E�]�w#1����fX�fn�*���v��[P���]j�c c���kFI�h��	�)EtKK��u������� �/*�/Ym��el�2/k.���.P'�H'f���*K���	Wŏ?[�������k��vғI��j�7��(��L5HM�,L���ݘ�Y�V�7^c���D4g�t5��>�y�zd���/��&���z��	@���2��A@���-3/zm\��d�@��P���d�>����,A7��"j�I���+E�ח�T���Z�5+'��[�Ț�%M�{���߭p���2~/����3��)"B����r�k[�u��N/or��*���|�ݥ��?d�Z�K�Lg	�8����6�g�g@[��rE��� �#�^�6�@�]��Q��teP��(�T_���r$e'q�č5\5F����N2���)�{釠�&�$�b�.B�E�d�65��;Oȼ��I#H�%r��ڰy�U{��>|co�~^�z��N� ��>}�Y�kQvD�d^� ۿ~�/���~uh?��i������wD�[#�h�ˋMR�糐�`��Q������e�~�,�_*�s�}m���'�$�y���X� �n��KC�z1�R	�_������;� &al�dvRb�5���A���c���
dd#FA�A0�+����/�T(OӠ?���X	���Ҁ%o��Y6�eV�����5�]���]��tl�X�:.������[pM*H���Ӎ�����N�tk��6���rp�̿�T.���6�x���9���k6{u7��ǡ*|i#Kr�G��Aæ��K=��yynl���h6*��#�p�VrT�Z�Ɉ*��`n��０԰�ɤ���Y01b�aY!�b-�c�����B���2V9"C�m�y��,�MP��˓ǌ�}壻��i��<}Y~i�9j�+޾`^T�g��g����EW���
�`|����P�p(���D���툭�Υ�Ug9��f�{D����㥺�w��v���xn�_y�N�$(\.RFNO���d@����t�}����Ȓe��ۮ�a���W�oPPЫ�/z�~�5H��X�"�UE�fC��  J~<#��UP5�q����y�Z��D�yF0s�����"(�c��$Z�(�8|{����:����� ��u��#�	�Zc@�J�v���7�8b���GzxE�N5�j�q�GD��;"@U�����W������oe���w�y�`J@0ȋ�� ���8Kz�\F�kR�.E6^��Ś��6f|�nc�e�ۛ����y�5@D���LÇaDa��ƍ�A�Gl﷤���U���N�_���rV?���r���@����F~Ɣ�e�K��"��ƞ��sO,*��J�Аhb����#�i��f$����rW�0����E����N
(�-֯���\[py�R����3R`_���6�xxˣ�њ���/���WN$gf��X�� C�t����_�z���qu�ݪӼ�c���P����R9�w�o7Jf��$�$����8e���u,�b
V�|� %��8E�'�AZ_8+�*��v�*o��ϒf�]�QA�T'K�P��w����JO��*��<dw �z*#������Π� ���KvUL��v��p�V�j6���D*��3�����w�m������=F�s$��ʱ�-pu�@ٛcMm���]�����trJ
��sWlN/vx�u��)f�3�r[�{W�N,׾f�v�"7�i6�j�{A��F?_�1\�ש=�w"n!otFg����p���Í��_�$�A<��ԅ�.�' �\��,']T�+#Uѻ5ɢ0�b:�� �����o�GŅ�T��v��u� �.��z���>j����Sd�՚:�e�v�WAś����NI#?<�?7���M�wH��j�cn���İZ5`�����aۂ��PO}Z�4T�a���6�I�w���^�NC�m�Pi���4S���i3�85:v��>v#;�s��^I|�2��Wg��H���/�������<T��,\᜻�q��\�M R���S�-t�L�g.I\Uy绱���w)ZL�v>B����D$q����ZĮ����90gԼfTq��k��������)y���B��@��xL��w�F��� 8	#.������$k#&����k��lP3�)�ڈ\�d<�����0��F�s6�����d���vʖZ�*1�ݷƏC���a�:|*muyO�L�zO}!����莂��(�=�g��i�����Yy?~�i�4s����$a��$������f�^%����r�m�A�u�zP�A�v�hm51��}=�MM�u�C�v���_)D}��v�B�rߩp;�RM��;.S�:��w����Y�+�Z�̺��[�w�F��Y�)`�h��`�P$��9�ܸDѼ9�K˼+*����XZhĪ���[Ggq�l��4�]���'7sT�]�ѿ  �8 ��@���=h%��RLxL�˸��K���贕�wL���`}�:=���'Q���a�����5��>c�.�z�8�!bd7���K��RRf�w�!>�$��R�眬�9"����Y7�IY�����[�mo�R�q�O���qZ�6�1md/�L@���SW��H��La��M.��Ჴa�vݻ̈́'�E@���&?��;q�T�&L�kp�B���:�5�x�|���ٌ<#˛>�����ٙ.S����[�!B��~1%O �����v$0g~�|O��5���$�!�xi�+S*cEY=��H�V���v3d���;��t�-c��$}����7ֻ=җ�a�p��p'��it)��8����{�)EE���/��63Xz>�]�h�4~����69.��G�ά �+���j�q ���Tr�*�\��&}GZ9N"��g6󔱣٭c����n�]?ρ�+G`���Z��K�ƭ?�Z�m�T4]L)Է6�ye���*[1/�_n�Dqox�.J:�[��h���D��%)
PQT��:���44���0���{��$���J1��%ѥ�T�S�L/�V����� �NY�Kv�s����:�W��{6P�W>�����dB�k�j6A^ճd"8g�C�t�h���J%�:��qMEc�c.u�%��r�2Vw��m��n�bAمX�:��g9'�r ��O�d���=(�\���y4�/�K�ꌌ�n�\W��A�Qe�v�G�����+@������l^�ww/���1�T�3�{L�d�Aʧ���$��l�-�Wc��T�/-�9�W�{�7P^B�Qv�>����zo��h\����{���`}�(���}=\���n��� \ɿ�Wd����*HW�w�y+�K�V���]�G��t��������������v�䫁�e}`�(�#�՛qa|�o-%�"���i@�D�o�ѿ�g￙K���&��MF�����4V �ti&�ٽ�J�m���V�!�~7B�$H�^��9���}#�L�A���`ձ�t���#�дf�����E�s� k�|`�m�!�Ljz�T���d�Lb���P~�;}�s)�g�o�kj������L���W�����ё�zňF�.�_���a���IR�����B}�Fy�0p�-� �5	@�A�]���
�^����M�D��(L��A��O/ā�#D����k%�ˢ= 4;�������n�(�.Z����Y�[�)�M�˺Rs�E>gK���j,�):Ϡ�ʕ�F�X|ҷtv&��>ֽ��x�h%���S��׏����܋=$g���=�����n��%��~�%�h�=	��r�sX�|p�<(Zsu�0��!^-����h��OZU؂�Y��6K���~�7~�s"=�o3�e#�FJ[c�^2�8�1�n�X� "T�L�%��8-t"���k<�������x�M�N���G����rV�űa��h��hg޲�/���\H�v��/�1�u���e��P�c��0��⻣aagO�ׂ���^�O#���Ay�y����;J��s��/��&� #J��(m��MJ~"����dUm*�@mha��-U������1�a�rz�L��I5!@�r �y�ɉ\a��l��n#�:|zߵ�"B�"*��U=�{����K��a��Fu~�2�Tml�j�~Q��Я��v����_U��Oۆ)`t��Xpf�U<����*G����1�$��Ln�v�5nTE�G���� �>(��.�	-8���h�1m��y䊖����Kt���=.��&���.+�z�Cd�Т��p$�>����V��x� �-��<U�|��/@�n�,�ݖ�W��o���/=g�%���hy�󶳧�"Mp�ꍇф]��!��^�梹N6
�|����M��5�o�ni1��=�g�mbPZvvTFiV����WO t�f��$�l9�I�XY��7���ޠ��5�lK?�˫ّ���~�9��V�����}.�(�ש���&ד��l�Stn�V0P`PG:P�����>�V틽�ۣ�����}1���6d��T��:�?�V�:����^�����r-�%\LT��J`�:��v_U��D��\�=�����.S�\V�#�\Z�<f�f�1����ԩ$�y������ �z@Z�NU�{Z@~'�?���tY��;�-ʏ������4Q���y}�IX���Wۆ�&����U��*��^�r��fV�����"�Opkw�BU��vo�\f���w�͵�����ޞ?Z�(�{p�ae;6��N�� B����97��S�_<��1��V��� ��C���×Bmu�822S����w�<��$g�T���g��*�9��>���mK1AZ����(�ޡ��_��[g��(�5� o�@������$ҡ6�A�ψQ*I&+�0r���Q�Яl�}q�}n#�Z=�e�Nq4����,��@�x�a��]�&+�]���h��u��^�v�z�P��o���H��{!w��P�q�I�rs�<���>��� �@�y�g��4Vt���zC�Fq3����Q��l݆̍�0y?�ډ��Qs��f+�ᔳ�tH�}��T���P��K�'�;�ks�{�#~�e�;�gT�p�WVW<E�Eg
)S��^�P�/�'b'v��o�G�;���+�"ك�B)&8����r~ӿ݂���6�!�Lc�?�%�4���B0��đ���	)G��lܚ�n��R��ͳa?]��ܫ\gjp��
�:�@��S�����v0�Q'�o��sȟs�uo�Ћ�G�@T�^�b��*���D
P���}�S�7q�}� �#_Q�>C.�c,]�}~ɷd�.x�* ��q � �o�qcNm����7?�gǦ�Kce�D���{�4�\�F��&;F���_��~_�Q�.���r&�	d��8q
�D���:���>����bB�N?��P�!��� t�?��W�q��*J����Sĳ9���Mb����d���j�[�ɱ��˱��pKg[��c�
g�!�Ѷ߀�B�@� e�Zu�Y���2&܅4l���t��9��M�l��2/ NU�w*��bD�NC�#�4��a�/�����"@(Ա_�5�c���2�����N悖�3���B�9��-՗]�4�P��\���R��{�S�<Mw �ت��H-��e��+cɬ�1M:��|��������=�6�Yp��}mrr4q�����E=L�Yr�L!h
U,�0"�"�%��5=��T��y�
���`����Vi�?@<���ϸ�Ρ ݹ��_\_W�ŭpp �4z��qc�$�V��{�/��zZ�9�F��C�g)r��^r&'|l���&�fg;��T����]�GJJZ|�)~)u �!|��p����H!�i*f���6v�uI�����GH^]z.��o����wMP�l�nq\}Y'�d�v��\�I�4���t�k�7L��Q�%��NޓtЯ�V���TO���#��P�a0�u�3XC�?�1�z�P�q&ZZq�� ���o�571|A��Pq|JM+��7|_CG�d%��ZW:��.��ȡ�\yu=0���7u�!OGx���פ�+�w�F�i����CB�z�8�ٱU"�k���a~A��Ўxa-��s�j�(��%hTu����v����H��X%��G~L9����U�*/��+����>�$�r7��b��"@�#�����	�L���k�7����,�A4xT���"H$K�<���r�y� k���r�1B��h�H����/R-R��[éݱgL�BtH��:|�+�fNG�嗾"܃AY�CĲ᫸HX@c�f�6,�"#�i2��ɂ���NF)|'t�^M�.ُ�,����B���4Э)ӎ��g�o�>@[�'y{-�K�!���:*�EgԷ�(g:��X/�>l����{A �8^R���bԗQK�1��^^��N&⽝_���\�\@�1˖,v�$�S5#\���R���0�}�<��\�TJ�����o���"�HkԞ����0rb���\Å�a7��2c���悔2������Fp%��Ϗ��1c3>/6,,��A҈�￷�"�F.t�P38N:h��`��ॿ��;����rTπ��=}Z;�h��p�q�v{}�r�{2��p�ҜU��w������, /�xqD��@a,�֓�w@��-0�<w��h�;��BК��Q<)q>EU9�r��%�E�;�pa�����>jo�Ǒ�ڣU6�FJ���V����'��8g�#�J���|�c�k'�]Dl�|=�7���3:�!QfU��#���^O��f,˩��A>���MI�b�v��ڑ���jxz|~��q��6`�G�˚=~㭙�����~��Kg;�&��.�{A��\��7*��n_;�	�Ϋ��Gwm��鯘���X��y�wa��P����.v��6�D��aX�QK��Ƹ��n2�j��`s2C�ޓ��O���e�*�ngֶ/�]�-�;��ot �h� �R*�c������*Ⳓ,�GV��=�¶0l3ih��dWG�Ð��V���y��#tV�Um\��	�Uh�0�3��?�jgFx��0h��J�$s����P6V�pkM^_� �a^a����P�CS�Y�q� x��~Z�$��4e@&�j���F5�2�����Z����U�'@	��� f(a#9 W�)�Dh���<'4��B�Z�b����CK��k-�O�pg�۞� &c6ȭ�Z���=u���)���s��O�~�=����?���['d��,�y�Z�t�:抣i'n�t�e���.� 9�uS�%�>-��Ce'y̮��8��B�A<���t;N��D�bL�4�����
��0��KU�w����[Y�W���A`��w�"�����T��_�+�\uX�8G��T�J$���b�~U�@yNc�%������Md���.��;�>�>�s�������w����,݊��[�0����2�d������չC�V�AM��������,O�Å���Me�^�>���*	*��-+iG�e��} S�(�]kh`0�����%@B�Z��]63����Qp`��
�a#=�)�*{צF��t�7/�Ѳ_�����b�I}mA+�{�h_�CɩP���m�:�YG�w������ŵV"�1��zA��a~��U�)��ߢ2��H��H�]��LV������0�V�����f�us�!���j���:�@^��,df��k0r�?���� ��p��r#[8�/m�s�X�VD�p�$	+���ԹY�?�c�&R����2m�o���Ƈ8�\o�ޗ��L�Җ��=t8�p��O�99D��k�	���o�^ӏ�t�>��e�����}�䦫R�}�?���_h �0C�~g��s�j3��`'�N�-�GD�g��V�a)�dj� ����0ᰴ!�#8a�������g�� ���H�\\�Pn���X�"�+ a�j��`uyuu��i����{-�d�)w�h�_=�+����5iK�y�"����ܑ��#�x��pr��W(��2�	T�Fx�:zf(6���V��ܫ�Ta(�G<Y�&�l�kc
�ѝ����y��D�n�����h#�t��Chճ���q���u������%�i'�	@5��!5�ڹT+g�+yⱟ���U���ӷP�7Uڒ|�MR����Wp��S\#TFIn퇿^�:�q�w�F���\��h���<��6�I�d0���;¦?�Хx��y�s��Ua���ay2<����%a_V%�tF7|Ә���t���(@�Y~2�8��%]���A\;��
�����/_��|�� X�D[-$A22�D�J��U��]�����"f��}S��(��6�$CSa<�d5gZG��_}fe�8�3��v�X/�
K�U��'Z�@(@{
�����_հ�	���<������ԭ�� �c�Qn�������|�ư`.���[���4���B�&������`���|"��oa1��$|�=�<��ִ��+�]ʥS#���YDP�bcC�܆�ˏ�� �l�BӶאF'�g#7F�[�+z��hJM��Xx��Wv����%��9X2|ٕhKp���+Q�q�e�xT�{��̡X���A���}y�M�UY�
���UMp�":Zuw��,z(٥���p��17��#�(�,�-����03,&���xx��
�����<�l��ё�3�{ٟJ����hd���ʯ�{d-xU}�ћm	�c{n��K��m��q���
�f�]�n� J�W_�P
��n�$����<L�ͱ�	�u�Hz^u;�C���	�/b����:�sCy�'��?h�'�Fy�� ����sQ��k)�qs�?�_?8}Op�Qt���I1Z�;HNIy�j �VO���94q��s��|5Sa�Ȍx�Ɔ��Q�>�q���Q��N(����������.z]h3d�R|����"铳%p����G�����8���0xG�����#ȃ�S��}y{ ��.؁?�M\�UƎ��!����a\�VA`�>4
��Ȇ+Y&��;�K��p��^��&�ggx��\e?�c�{H*�ۮ�أ:ۈʧ��1W��a{ۜ���:{h�/V'�� �:���:�x�$�ȟ��X΢�~3�T\��}�xϜ�`!w�����u$�+山����?i���Ok�q!c�����E�஡'����=��=t@�O�b���&%Y4Z-j�F>�E��ac##@�7l��2p*����T�CE����W/-bq��d����פq����V���&]|���/�@eL��E���n�J��2���#]U�hE`қ�ͷ�ē�N�"JF��<���P���(��$tkf�rf]�>B�3ag��t����4@��qxk�@�:*
ܼGx�צ&�$�"�S��ֵ��2]��9!�����A�`���[�pa�H�:/��<�$*&�6���y0_k��
�=3�u�w�f���i_[���Hw���:F"���|��3�C�c�X��pg�ecA���+��0�D�`х����X���O��rR�)*�<�|��S�5�P�ְĜ�v��ʕ�GJ��ltΙ�,H��UFO��(��tǬ�5<����++��H�C�T"srh���m9�w�� 5�;��Ї��h�k���#�Sx �FE�ҭ퓾���z�u�WD$�����e���%,88 x�>�~����	�V�!L~�����n7��-��I���zX�M3Z����r�������ut��5������s�j����#a�B�?Ĺ�m�6�QF?%���h�⚠]�W�������u��0>���iz?.Uᗉ���.�+�wJ(�@�}�����u�2�h��6�	�k����p6ʹ^��J���.kon��qk~`�>�G�A
��ƽ�ko�iw�nw��8��]y|	W�p3��ڝd``�^��L[��;��@��&N�/C_el��te���7�|H��ż�=q�14��Fy�{�Ju�����2�5[�W�9Y�}��&��E����L2w�m@�-��RM5A�._�PSR�<LB����(��I�.�8�$���h�U�d%� ����6Y����P���Q��J�;:�:�W�DF�%33~2!e����xSh����M�%�B���5���x��"^�O�+g5_B�M�S1%���9�d�Vv~�/b��C,����ET�b��� �`�9,7�L�\$"�2WʡNZ���I�ᡅ���T��GE�R;�t����a���T�f�H%����#�`s�Y���1|n`j�L:[��vx�7��ad��V�$�r?��mǙw�^���:���	DЁ"Lr�M9��l>r�uO�(U���cv&�c}?C���+&YP�(�ѵC�e�HbH�����J��M��l,|S�&�,M��v�o1�?;���0�{cMU�����@υĒ=0:f2뺗bV�?��������ku��Y�������߸�ʢ����9�6����t̸*��a:�<E���dg����`�IhCk�	ӊ���`��-R&�p&<S���'�S4�ɍ������F8��M��!{FO)2��n�wq�.W�;U���qUI�i�_��3E��Y*o�����h��j5�N'�;�5��4 �:9rB<���,^4,�}hI")-�*Yrj����1p��,���B��b�K�@�g}��.a^R��^��F5%��d���dk-W���B6 �NH��Z��I�,Y�i3�f�Z�u���ߟ�;�K�q}j��$�Y�]�7�]��nN�Ex2RP���Y����	\��[D�9��L��f!^��aY�������K{�ԥ���}����x�{�d�Mt�(�v�@��e#l&<GKDewv�.����60��%��,�F歺�t�'.�}�Ig*�-ג��&�A�w��櫓7���#��]9���'���r.o�5r�}W��z`� Oa��|3	H�6&v�5�ᴼ.(��»᥃��b�����7�@����vPQ��C\ȏ�`�����J�BL�ƺ�p��[
��M���|�Q�òz,m��i�%���v�P�����F���M�H��E5�C��nS���E�W�?�[Մ���{=�n���Zބf[�Z�1б1�"f|��������V</Go[:�^eS��]���*�l�4��&���k
Q˧&R�81B��NX?Y�r�Ϋ��V�F��Oϴ�IB�+{���͜aq�������X-�|�Yf��FR5�|�{�	��O���i#��g��;eB<sV�**G6�/6�
�pf�3��{�
w�·��o�"�Q;���v;�XӂS�x�S���W>��pn'%�@�"���+�n?�����eo�: ;�� ��Hi�~]0'|�`���B���h����@[z{��9��'�k3�֛#�td�&��&?~a;��]�\�zpE:0
��CP�y�fɂU�6A�o�?�7�7+&޷N�*�وƦʝ�i~�l�,��P&k�t�K��D٭�����z !��8�Bʉ�HQ����F�������e���U�3.�G����y��ˬ��Q~)���Z��?*oؚ�z��|�09�{w�T���������U=�Z�����	���	@@���ú��F=�(�I�W��1" ���X�0Q�Q9��i�0����;�RD�����?N�I'���z0a�Kk�0� �OD�~���Ta�M�1O�!��cd&F,��P������#���5���~���qk�����Vg<���<���0�h�e��ӗ���zo����F�Jc���N��W��74��c�Sg���R2��Z�j?ػ��p���9z�6}�ҥDb�]�u,�2x��Yf�+�z�m3��D�2>q�!���wV�Z�X���:m�,�"��P����й��͗PF�K���Է"%�Y.�
�6�P�B�����@|�xM�J��'���0"�VWs=��?���,w���2(*+ϵ���֓۶�I�d�1ҭ����׭�p�\zz����+���9���Ֆ�O�!m�h�G9�p�5P�xT����`$��o2�\�MJrR|u�H2��o����C>'��]�΍K5�\-�̠[�<��0�Y<�Δ����
ysd���ji�!���4��rҕ��K�,/���U�g�	?�L�҅�x�}%Q0�y��\�B!! �`D�6���M����wTN]DxM����n����}�"`�`2�v������X*SGǏS�ܙ��HL�#�a=T�z�#������I&u�����]����ޘ�
�?�����ի��bS6�#ӗ���)vAc�vߦ;N�Υk�.�_���h�U[苭y�h�]�Xq�렟����C���&,�۟�os=� �� ( �{�}�9��Y��� MZ�
o��Ԧ�j��ed��2S\�"f
�(4� �ܰ( �ӻO� ƕh�c<��*~�+��}�/RB�	#������n���{!m!tKxv'u����6��������;�]�u ��#X붼[u@}�_�⩁�:.��?�9Ŗϗ���;�~��pzl�[�u���!i�D�T���=K;mg�X��x-)��`<�څ�x�1�Q�	�1�{&u�H�����7G�9qy <``���\χ]4y�3z*�RG�c�J�XXp1ғ��!�ݲu4�M �?�/�qF߁�ˁ���?�ы&1܃�$1��@� �!���5�n��+}Z��v_$ 0~i�-b��θ�3��gV��~�������-�S�+z�	X4��CR�/8Qb��K�K�xUNإ���=�� PU�Yz�D���� �a�3����ǔ* �4��@���"�7Xd�Q�(�K�R���W����G�O�q� �aY�s�/��^D��t ���{ �����W
D8*������p�k#wwA��cb�6I�tx�`S���8m#���5PD��K	�g�DJ$go�z��+9�{"�BÄ���0��;�,>ļ����[?��� j.�� ���	ڋ.PW�`bĨ-�x4��j:�؇�4�Of��W"�b������Y�������D ���/r���g�G�>ɿ倿��qo����������!wח��O����t�������'��x|H�=;p�{k��v�HeI�{$;�o��`X�|m<���ߥ��l�<u?�t�^4��=�~3\¬u:�����W�Ҥ�޿3�p�j�>�u�oϿ�Jh�f�ʒ|�,N�ܿ���/TK��������-�)��>TK��f�#ѕI�X�KK2>�21ʝ�e(z�E�Ow�RZ*� qeb�X�� ۊ(����.��b���St���"�h{~,���^��/��]�Z}𶀑VZX^B���B]ő�v�o�j���~�����v@V�_�%H϶���n���|l����fC�}R��Y�a;�ϔx�Y� ���h��?�6,���[h�`��V
#�2�㔵y����~;IX�]�22\h��$FpD���xz˰6��k8���݊�;)
(�]��B�J��w�"��C�Bp��%��>߿�G�s��^k�^{�Ӫz�|L)�u<v�*f��wg��$��d?u�B�d�іٗ��C/prr�X2!/CR)q�i�����Nf3�偲��&�9Շr�4̜�h0w�kc��p�����4�9L�y��D�1RD}'��]�;?�.*�{Q�q$�����[p��ѿg��=��s�lנ##���n��;�;R%����[���~�F�M�����%ݷ0e6^��y�8O-1/r��Jܧ�(��O;p���B"�
��٫�.�y���L���� ����e|��7C�필ӈ����9>��W�3�� ��FhV!�&�f.
�ƕ��W�s�	]0x \�å�Sa��b�e��inS��-�Y��$�Q�)�(UMVl��j�o+���TGן+Ƙ����3�8I���m�w�-9�K�{�S��ŗ��N���I޼�C�u�{
:���{:>G9C��o�q�2C������r����Ҍ��W��3 �w��-Ї��i���t�"��X��ķ�'E3$�Ȍ~Sx
;���8���`ec�q�Pkn�d�����񊥪D�i�] �9����!8��5�I��͞�]��wc$TT�\�2����D'5�b$�ߪ`6�`s��"�J��8���-pI�o�J�H�ߏ"���������+1��)Kq��m�Jl�f�L�:��1���5)qZy�Ej�G�6{!���ơ�xs|��s���M�gg��ͩ��X�C�����N�������nuEt��i��J��9��F�Б�>t�_�Vc��RK��U�����o����SP�W):~t'��-ϗk{������.}���M	��a�oR��$xdC# ��n"�&�|L��8�@���Us*��ñ��#�g�=`�x�"��{��]�t�Fm,}�U@��>G��P�rꄴ�$�l*j�8�g��
Sj��%?��獁�Hy/7۾�[�ô��,�U޹ś_��<���p!}pz:��o�4m�����u������M|�T���D��m�����'_iP���(�B%��`'�d���[2�f)be�Y@�ef���D@�Qw7x8�i������O��`S���"������9����:	��$zS��p��=B� �.�,+*��7  �ܮ��>�c�*&(�*F��4�"ΌMwvo}ixkn����T}C��
�F`�5hk�p{ ��0�����: �@ʗS[X��uG���[����h��;;�}�6+�����3s��<�|�,�/��t��bu�����"������I!���T�Z�������xo�)��~�9U�.�ke��_�f��t)��'���'��3ة��߆Y_Ts2K�#��C��k���C�-{q�������"��L��{z����+߶E^�P�<IS��;A��A���{�����������K���P5�6yDڵ�S&�PF�q�_+`6Z�O���W�������tG��<�03/\̰:���Z"d_�M�?s>c�m�]���dx��o�5L�]I�sQ|	��,_|:AC͕������6H��Y�*�5��?�V��h+a�4�V�'n�}��֔�M���u৷A'e_ot7�kN�����me2);5�X�i�3,m&Ry�9�qE�kG��. Di+�-A�m��=Q&�5�a9E��.8�'�Y� �k�だ���0[h��>�n� H}��=��0�8i����?��ǌ�d����"9%��ز2vɳDwW��㩗�)��/3-�uhp��ϷTw�q2�y�H�V�i�����u�����_#���o�&/O�+����W�ؖ6#��n
 W��>	<��)(''QZ*P̐M��KH���K�|��$�A�-*�"�\Pxd�'�����h���7�T����_Q9�ߡ���,o�V Z�r�w|aNw.��b��d�߂<G{lG�{Zqy�2X�껶r�8s YXY�ż�j��7��ǽ��D��/���e�Xۇ�� W�6>��/��a��.��a�B�*E0�v1�H�3Q�x�R�0�'iʥ�dr�S9�	ǧ�}�/kp����ꣀҢ}�h�O}��h���5O����m�ď|���ُ�+���e���9xY�k�#��#�'����nS���N^��L�����)eY�Y7MYmq.̷Ll���{Q0kױ��(�T�*��5  �e��̕�I��1�v�jzuO-��G�<��	�:�u�S�;T�ЮZ�'#�� �R� �6���5X"3'4�3�� 8+r����+ǓT�8��sL�~����6ߟ�%���}9���|G,������?�D�͢;���S���bM��C�i;E5�|���`Jج6+�%:5��o�z�V{f
Ǝ��_�)*J4>��q��3�ʻR�I#} 	뷨�3,B�(��_��Ti��p��|���W�eD�߁���\���Z�O��H�T�*o��?o�<o{/�D��ru{˘1>�|�~�՞ 7�ϼzx��Rҷ���8���F�I�:�O�oe�Rh'n|r8��.�F�H��7�h�?S�����y�
��T,�P뻑lp;]JW�;D�5�U���KFzkL�n�����U���#J�*��V.�O�2�x��-l�������j�o�P�����2��;%@��Ija���o��?0"�ҏ���lCO_����g��_�1�>虝گ�I~�����Dl<���bD�ia.�O�ˏTRk(�OODb��S�,��@�`�Vi�#����kJK��I�DօD���Yt@�l/����� Q�Ճ2O$����
�c��ST;�G��J��?/ 2�̡ǝ*p�̮m1�����c�处�:O��Sq���7$��E���HD����v��Gܼo��"��r�f,�jqu.����}�ؖB��U��+w���g��ᩮ����� rҚe�0� V
��#���e�W3lҩ�4D}���$.ˡB� L��K�8�_�*�?��Z�@� s�WFt#ƌ&R"L��MQ���lݾ��O�M�H�|�]���w� :��]����p�۰ge�u��~=�Ԅ��&�@E�_���������VO����ʬ7(���wpw�����a����'�ܻ�Û�Oo-^N`d��QH�$b&�����Qd�]���K���i�?��}�x�r�'b$���	�Nb!w�W�#��>a�+�����t64:�o�
@O��y�\�s7�}ɖ����:�g���9���:����x����6��g����uSi7��[�~V�'�����l��MhSsN�����+t�H�H�reL�ز�iF�$��e� ܱH�̱�u�%��F�"9�I�E�g�~��8!����� X��7�!zBָA��u�b{:Y��^�qrJ��e����� ���%��.����N���[��'�÷ZS-���7��"�M�����v_�㓑,�[%�7/{$��w�(r'�*V'�y��_���Ƿ����{�Q��K-���\�/5|�K�!���Oy���9>0���hp����v��E	���9ү�i�g�8�e,��&�&��i>q5��$��\0��腙=m������zQw�j��"1�IR�vGY���>�}B"��b���?�"=zM��Ӓ��r�3.�ȴ��<[���B�8]-��*1�ZY=G��+пF����&a���R�f�����o�*���aB�/d��F1���j�z峌�twgtS�^�<P�݆������l|^o8O�G�]d��p7��d@,��	�Ɐ�����F�ʾҹQ#A��KW��հP.��R��򷍌4�MYz�y��TA'2�l0=�-.�/0�K�h������[n���o�-��IA����[�ǖ�c�-�~�� ��x��)�J]���8�R�J�"��hv��0�ۊ4h�b��}�O���0����3>�K�O0��1|��;�Yb���il�F��������C|P��{��,"t�*r�&��"�y��8_����[O�B�d�~��4�m]�>�����<8&|��%����F���L�@6x|�
N��Ic<����UV{�hE�D F��S����G:G���X����aiA�	8#�6M�]�����Ab}�p$���l(���dNl��I����8��;D�<�&��"�g�a�L���%f��|�m�1��hlHQ^�q|��
w[��%���x+yŲn 8�.l{�pyz~���k����[L=��7v�mga^���~����cYo��T��.��?(��M:�K6=8���e���@Ba����m�y�����@6M�����]ch�e��7�鵹�(�nG��G�vs7��_F�n�C��|�:#��D��N�S�Hy�/��n=6��ϰQ,;e��6�Y�w�`QP#ޘ�`�i���Z���/,%�_���HlCi�>�?0�&4>����ƈ��%`��Y��t^i2_�6q{���������k=F���K�����q�y:HMf'�%n�"��
��!�U@ ��s�g�ǲwbC~"E�����O�O<��B(2��"�)��:k �fB:ju�;���-J[{���=&f���D �I��yEҴ�r�~��o�俰�M	 LI?:�8V��LI^b���  �9�(�g�r����MuU���u�/�l<�cb�k�~v6����*�2Q*�mСνg�����w������Ԗ���^�I����bL����i�bΊx���۱�v=��r��~����f;��s�0U8���V4�c��u�9  ��7L��
<O�=���8��?����+� R>V_���`m?۶�jG��6lq���+j9,��0��7�[;�&|+������C��F[�#�<	�.�hA���Td�#����b��l7{��d�.!�I����n�&���	:<YC�y�K�f��ԗ�4�R��G��p�c�g^?m\e��4�$w�SWՖOM�&�<R�k�o�f��i�/�HLR �p�|U$�꿷b7�@j�`�Bqf��A�j����}�7t/5�7�xu�h'��n����<��5�D�N\z��.�{��Q�aS���Ӿ�O8�~�
����'H�9��/`���u�+2�꟎"Z��*L��3��Ol�_�8�"9p񦋳���'"��N �!-j �r1N5QQڅ5��=�N>���ӌ�Gk�J ��
y��#�G�\ ���{�A�k�;>y�Y�?=Z}��>����<\Y���V�O�u�5�r��KF��5�W�T�O���3J�[%2����h��gY��z�;>z���W��&�D�j��yO�H�Ey�XL%�=�i|�����]|�3F�w�z�Tr�z�1��ۧV��d:�N�E�Iǽ��-n$��K�P4�� ��;rziL�U�J�}&�@�+�a�q�Sѿh��=�&�
�ox̍�%PbfM�2�7����As��L�v6(	3� �1�2�)�<( Z��J.�|/�U�ҏw���;�;�t*���~j�G���g�n���LQQ4�}!!�c�t"+�a	��X.z>%�����gu�3���Ԙ��}�oP&*lV��X�s��K����	���A&,i��j�o9Bd���4=������:ZE8�4� {�z���Y�����'����ܯ���L>Ԓ�W���S��k��s����D���l	��ݧ���ICvC�����S�3:WGX`��f��K(�+h�L��=O�*�֮�t����e2�alFi�p���Ȉiu��x��N�?>b
G<�3��oz	xm|��5R`\PXb�D�A�;��D���+�[{�޾?_��n'�͎��!6�_�f7�{�/;(;v��S���q���d�U��(d0e���M/W(���/�I��9�/
7`��o���Ԕz�����R#	Q����7I�����+��G��u�ko�ਹ�S.�x�t�7R7B�s�{�d�R��㾔߾T��c:��;�?��L2չ�
=8���m:�]X���nr��{'�˜ZdT�܈.s׋�!8p	�}�+�.�-����5�k�l�u�yxX�N�����zs"ٱ�9�xGݸ0�tb�U�b�5`Ob�IG QV�J�2{'73#�O������	&5�	���õ���?/�>�3�U�Zl��""���H�aܚ/ �`^Mo��|�TT�e��J��є`C����������!�[�
��;'&���<}�Z�}I�?r���MSF��Q7لw��"PLap�.I�K
3�&Ǽ�]WrjS�B�̎�Gƈ��5{ү�����W��8t�Ө���E��W5��qmq�^�2��@�~�_�CQ;N�N�:�wU�oJ�5���
�g{�NaV?�di��o�x����-a`���!L����� 'úO��Z|��4�i*����Q�f��������ͯ�����3h!Y!�n�価�`�T��G:r8)3P��77�T[0hM-�~��!�� G<��&�4��t�9ݧ.��7��딚܆��0>��wXdP�!k'��ֻ���
Y�]/���Z�,�p�Fk`��JF!�x�",��[cz�V	��0�Pv�ߪX��<��?Y��-�|��FH�}ʅ
0w"� f�P�w�w�=aȘg�\�	�}��`J����ׯ4!&������&w����_�`$������:��4G�}�W�5�'�~`�� �l� $�����4�}���,�h�e�������-�/E��N&BO��)�d�j1��G��ڵ1p�K>�BQ��C��I����F�^3�Q����ڄ �lU�F��X�Y�� ��I�~Z�� `n�z���ӄ���PZ�\�
��z7_�u=L���ӬU���#���i�A�"����c�q ���K����G+���Ujv���	i�������j���.o �M���#�����[��ۏ�G�P��OV�GJ�B��l@�����&g>oNy�I�*�	�N�u&��ud����Y#�jTQ��D��y�>(�X��0oG!����H�>[�� PW]�o�n���Z�
۸zܑ��}���'��J���v��\�$�/ZD�����j�X�ґ��8�m��/RQ�GȲI��V9�l���`ؠB�0][5/edtoX����2����s���	o'���l{������oyl���F�R�N'}�-뵮;���8�'�õ�Ȓ������}�0F���ֽ8r���o_��3^>3g��zl�Y��)��k�Ax˝Տ���ь-�K�(�B�lVv"O�a_}�3�w��v���;�ЈW����������+[�wI�l��6�������l^�.8���'����&!~��n�+�<9��X�+���ߑӀ�n��w��9& nQ���OU[Mě��5@V]y,�p5�k�<�_�Fd�|�o���>�	�1�����������0�}[/Z$�c�'�܀��c �R�Q|FV��ŧ�"y\��P����x�	��FT#��o�R����5GފfǪ�>cGo��6��I�����kBُS02y|ԏ##�d��\c9�zk4�)6�|�f'g{����Uy���ѿ������k�u\6��h}�K+�'5����ny�d��+�j�UIA2������=>� έ������D�V>a���}#�dR��2?�I���j�К|�$�xn���޽!s��C�r5xl���|���1-u�4i"�B��������Pm�n��^����\��/F.@ ><)�	�,���rQ�+�38!5t�p?�Oz�t�b L� >�~���~,^��T��X9����ى�8H�]�*�$�y���A%pѮ����+�OOr�j
��Ta"�&S@IF�/!��j8�4��T���QvCqC��O  (M,f2�g!�,����)֮
��.�Q	��׬���B�	��6n�.i��87"�ɼ�{��;�'��I�3����a���c�V\Ɋ
���Wx4h�n:%+�2O�A�0�!7��Kl�步����Ĵ�+;��xs�!S̖hhie'Q|5�!����b��M#�l)�6c5�]�'|IV�B�h�} �7_*����/o�25̌���E�W�Y��s�GX�� ��<#щ���xy�m�g�]Q%f !��ޤ����Nj��u��H0[�1]�/_�f���6��]��|������!�E���*�*��B�A�@���Q9d�3�t-	���jdHJ��A��zQ&L#7]�{o�@o�%e�Ҷ�~L������SC��vEl�LQx$q�N��zo���7�;n2�GP�����~�z�U�z�}��0-�1Υڂ(�I��Z1�Rd�f��5��(k^|I^0��� n�)O�N�oS�&��4!Ҝ���Iu0��[�o�1O�#
h|���.���:�x��l	�L+ѝ`��d�����*H(~1! F��|G3%ǒ(�\�1t�m~D���A���GJ~Ye�J���D�U�C���أ�n�)^���e��M�o�Hq��{ ���$����'X&-;�(+��E=A�ڀs��S�ll[�*���x$�Z_��k:���WQ�-(����#z�1X�DRk.!|�������\g��@���f��$~��W�k�dte�-i��!��L�����!(�6�j&���MO��P�~L��kdG���NdRcp�zF�^!_�#ᷠm�7�2��ѫT��=��$��앦Fm)�7�%Q��}���w^��Mׯ�V�7p�*�0���Z�u��(��+y׿���yS��#�Ʒ��ᅢXs�0 �m��ih�/`N��eƉ9 |�$�[� �I�dô;�q�2�Z�|�`�]C�tB2�%��&/rPD�4�Y3�K`.�Z:�8vK�`��6[�"�1�#j�o(�N�,��&���s!��� ��d:�nIz��y+W�,��FN5V�Mh���s�����bm�������2�i~����_-����_>���w�䉱jM�:�m�K8�%!���WsIZh�h��ps�Z| ������n��L��?�v��L�ľ�"�$���]Mޘt�2�R��I�%�g����Z���b�������g��A�F/5�Z�Ga�{��
�B��jL��x�ㆍ�=��	����,��q-�)��}�&�7�&d�D[�3�>Bb3�D��%�x�{5}]%�Q�O:��?}�$[���vl�X��7�1��Շ�D��)^)T�㾯4� ���S�Z�=�{���X�x�3����5c���C�4�H=��s�Q��sa�X�9�,L!
PBE\�d4U'����s����Y�p�5Q�� /��>����כvXp�Ł+cD6�;w�zjמ��Ͽ������w(}��۳z�c���c�p-��r����Y��<NL�K����X�N�=y�W�������"��~���0�*���m����ێmy�>����S$l7���oE�~�	:v�0�{y���3���� \��oj���Ѵ����V��}����տ�!�yY��	OJ;o@�ٝ�t�P���o�&oYݸ��o�*=���c,L4q���Qz�1��	Q��jZ�'LkOV��@:6�?l�6�F9��5�
�����b<��v�gԙ�F�6'@����Q���ljM�����?����L�)���N�5�z��n$֐tˤ�!F���mE���2�Rs�vS?�"?L�R����7_f{�DDR�|l$$��pl²�]ICK�m�$���tZ� ?�xt{y�E<+�|�[���,�qy���z������~K��J��4ZE��~�&�xcT��.���#^^Wv`D�QTQ) ��K'H֏����9�2�ϙ0�=���p����dR�\���G&���^JD�7@F ����Ǟ.`%R�����ށ����TN�>�n����{P��͌c	�>�E�m9�15����jz���Е��Vy]z�y$��aw���t�~� ��c߂��M������U�9͟5F��x=k&�4~�3kWpL��Ol���\/����gg�;�g�-{���1��7�?p�A���#���qU1
ݧ]�X�����G>��&����Z���='��C��J�%�rc����B|&x#�����v��xR#|!�25�ֶ\��f��ψ�~I�5�ѡ��`J���s��S@�D1��M��9�݆�2
�Ʉ��G]����Z��Z�:�7J�"W��-X��ʼ4�Ub�{�M���w����׼��#='�J�n>9�/4��1�$�x�6[��C�	{�C�k`4�s�#�J>�'u�}Ts�<=F��;h��i�&�s4���{WSo|�(�Y�[��B*�-��֏5��#��	��l����r��F!���+���F��+ }"��m6���Ó�c�(���R����<K�fv^��h6��J�����clb�"Fu�&�*����(�?�?�w�/�K�On�o�D��,mV'`K��9�2�À���԰=��RĤx9�34��'����K����|��ھ��.��Ľ��W�q�:e����	����Ό�$]�A��]@at?a(��̧gYρp�_�����إ(�X����#����)��� 1���-/�"x���gdc�����U����_�o��Bss�M|N;o��f�ݮE���pA�"�{�x̟�f?]g%K�M�{�N@�D���fq��r����F�#?�
\b{�P\����^ �y�Q��n����.�S���׫ժJ��K�ϰ(�JRX�nOV��p��w�D�^�Ej��Ƣ\�HS�G�'WN|�d�I�z`S4��{ �}�߬l9�+�g��ג& y$S��ˌ������g������C//�������9�j��l�.r���Wb�^����(��aEM��W�)�/Ϣc�Α�iGw�Vi;V�:A�H������D3�n�9/���VsE����˚0m���M����+T���d.3��=���WqN��Ȣ���-��~ �9�Rm ��g;���΁�R��6�Z{�%z��l���अĦ#��Q�֡T��0�+��ðQ+�ڴ�3���5gꩴ�΃p����q\��7\DYi_s��D%��4Hi7b~X��CL���P���_L����i�y��&�U7,s��X=�1d9�,����B��~'��߯�y=Or����gǬ�/j3A�NfZ����t�M�X�G�G ^�פ~Є�Md-�v*$���w6`�/����Ǩ�M���{M�3R(��n'�����u�����̩�z��D�n�	��Ď\]���΄CN8`���,��ǽ�f>M�.Y[�V~5���=ʉ�r��E�-����1>F�2�n脲8���p^��I��wo	�PvI)����Z��4��'\f���R�*��J8�1�k�K�uޣʠ�̩=��mZ6��T�\=���#9��NBbg{����G��D��}�%3>�ˑ�'����]�ꑿXo�v�H�p/�Y�_®4�h�+FSt��_�2�؁��6����*|6���`	�yk�㜪�v|5���T��6H��"|�P�5��{+�D��ѴC�[.���ǹ�U��i�3"T��Л�@�}����e��4
��4�A&K��	�S1\�g�d�@S�$�?�Z$|�	�"%x:��D�t��=8Hj����e?[�[�yu5���@k�Ņ%i� �,�wʏ�ӛ��B0|^r���+��3CKρ�NE;��z�������������P&���/��$A*a�������e�G�eP���
��O6��Q��]gӋ]�����1B ��`[E�&)m�Bj��B1�6Y� _[�R�%`�R���ڏ+�A��҄N �%���WX/u�U�O|�>�D��W��P���t�V%mn�T��=i�3�nJ�+4Ŵg�2;R�?oN��=�"I-�nzÐ1k��aa����?%�]���'61?��ѳ��א��.�^f�x7����L�z�ю�f!�����%��b6��x!�����S����w�����M"�B��ִ�K�ΰ���6B�5�M���.���5D��"ݸ/����Q�V�_a�,��$)�K�Gd6~�2�kRd��Џ�K��Z4�\ئ%����[=���J��ٗ�x(�`K,�}c��3����++����?�|QX�W '�w;�/1���%o��>���w0g��}&٥��a���;�M��ռ���c��I�ڼ7���_*\�p�U�A1�X�X�͟�����y�E�!ͥ��}���1��{�cF;*��<����ʨn��[4G���s�U�{��9��n�<�����abvϼ��}��ɳ�����?NOd>�.Ҙȵ���R�M�]g'�+��q9��r��[� ���|8���݆6jU�<L��C�O0_��H�V=�?�?K�4kF�m�5�F��'���&'��iBY���o�3�;;�u�Z�ژf����;�͒1�f�������;��R�Z�Y��}� ����Ͳ#�A-���嗌r�:���rVT�J�Mb�Tg'o��;e��,��=��W��X�����ǟ�oL0�ʼ.-]��گA�G4���������D	��J !�:j$KV&���p<:��8��{�JVAb������yN�I�AW��.]�z���`����ꣿ��<��x��؁�J��0�|���_�SG�g�C6x}}M�I��i�3�ϱ����әK�a�χ�|�ه��	�/� ���Gf�W�{�sx�糊�r|��\�ڀ��'s�F����"x�z���y���y�����4�O�3
mf�;?�������ۧz�-�]�_�#Q�n~�ں�����Tzޱ���BN�ͩ�S��?g|w��[}}�Si�R���,��7a�BA��n#ɶ02���_�S�35ܠ�򚟏�G��M%��1�NX
�U�`�!��SC ��\Tx#1�]:� L�	���'�tO|�����V������l���!@���M��S[=�TR������A����"�`M����O����\L2��h�P�.3��n�zw2]�����3O��;GZ�ІS�Ǣw�7�CT���P���}[��ֿۗ��#�6d�ĭc���
0�r/�������;��ZK��OaQ&\�;B�֪��ټڍ�G��?e�"�3�g\��IN�<'z߲���m�<�xM�ץE�/�j2GLt+��^%|wd���2h��^4G�9�B�����ɥ*��9��ۭ�˷�BQ�!�2�F]��?�O}#�A�֎�%o���≦�C#d��q"`��+���^t����f��YLX �����'�<O������;������_5�!vy� ��#ոG����V��� JߑqD�݊���^R��	.�����4R��V^���y!������;w�*���z�&?�s dY��,��n�*��o�W�O1�����E[�`����j��6�&ƫ��C�nY)!V��zDV��u	���.��9���-sV��(��?Ƥ3,�o� `�x2�P�Ki<`����E�]��-�\
�Qk���&��s�/F���&$�M��'���w��eV!@�l��b(�2O�.]�6p9��dc�W����u��9�
=ū�it��8ĝ�!3]�ب�̹R:.�������V+t��-+]���E���ʪ��N��{PV���@�^�%\�m0w^sn�$V�N�|I�7J�s��´|o���Â����^�>��f��-���3�7���%�.}FϿr2g^����bz�2��� ��6��DDoW=��s��c����������Y#��
�G�3@/Ϸ�O���+?M�e֩6,�!�0�S��G"������T��+���[I/Bc_�ne��#3�����Q3&�f�H�dk|��F4�އ_�,YN�w%���V-3�;�B�W��R5�eECjw�&¤���N}z�mGJfT����̿�(ޙ:ı[�
' x^8���H22"%����ˁ����wy�75�F+#����BY���3+3.*Yt$EYB�1����v�+�W���I�6J�9E/�p�!�'a\����a��A/n��u	������q�/1�ӄB���[�,R����8�~T�$�=�!O;�
�\��-�M+LK��I�����g}�[��R3h����x���j�$#dIͽ�-Bų\�g����n����'x�=udX>�f�3��:J�����[�uc������c�p��⓹�#���[9&3�W�<���&R�5t��̬��t���
���徚��:}��A����@�C�;U�2�Ђ��0����L*0Fϯ��Aq�T�y�td� �,�eQ#���[|(��L�d+I�[���
܆��ITd͋��D�Gĸ͋�����gZ���M����8������/��f��n�����v�[��v�w�|����
:�(���YymO�D�#�ܦs0�����~�s8O���u�~e�q�1����Ru����*~�Z
��[����4��bc����<f頙�P�Ȑ�C����,�``�(G*5���>�[j`� ���O�ái�=!3�e�%�Ж�:O6��-�3��!��g�����Gi狏�09�¶���~_N
9�\-��9��A ��1��{1P����	iM7�<1U3 ���KB���[�.8��4n%x�_]yT��'�i���7^u�ҿ��!�4`�U�K�38!�W7/�䷪Ӟ��]���V�p���K[=ـo�S�x�{7�[��	^C�{���:����gE�P�g��!��{�У����:����U� �������'`�<~�{�9��E�P��0�~+RX���ʣ���[�AxQL�����8f�ɷ�mؐ��j�4��
�eٴ�l�qW�5 �Ʈ��t��L*L����u�%C��Rm���Ҿ8���������U&�\NU�B�D��L��P}�4L�i7r���S�R��MJ�]s���q��z���}-�|���	�������p2_ռ�A�[]EdQa�l$�mngKu�]ns�w["���~Q�=�-���0|�|���Q��L��H�M~|�jH�谍W�(5�M���U(�X�ƐA���U��0�-���r��ve��Ւ�aMo���u�U07����Y��P��~9�ߍ� �>�`t;A��&� ����β���O@8�b�H�l��b�F~��J��~��ō�������Q&釙D��k�ӗT����s8~�UDT�`Te�&Q�.�ܼH��-}��z���kp3�����0.:��9�2sA�O]�}T�y�H:�� 眄I�v|c��H�tլg�#D�TM��u�j%�o�[�6��	��Ž=1;M�!˸+��"y��F��-j��*�#k��dK&[��%��$L\��5�"Ԙx,��H�ԋ�:'?8�v�'�
�3�7yNI5�=�y\�RcYIu�y�����+t_�;�pF�y��р�c��$NZ�^��`�j� ���������S�ݙ�o��ܸ����ά,�e�tt�l�����v��:�$y䲏�\�]� {����$-U��#���K���]�	��*�`�4��̘�ALS�'\��*�gӵH=�¸ �R��T.i�Ky�o���U�gE����[�����bEoD���fM�^�:���zķ��X��i^��_'�??s$-A}��UbA5��sZ�	n���M��8�?ڿ�	���)�����伢�<�4�~�?%n�m�A�Ռ���mIp"{��?_iX��
�9�T�WP?��l�՟6��,��"�B�X�$2ޚ)�rX��K��
9b�8�4*��7�ޯ��aYݠl0'/���Z�&;��Q�q84��ؠFԡ�2��%�7c���PZ�LQ<o�r�?� K�� �|0U�������lu^U(e?x�ժJ�A#Jd��>�<I<A������I_����1�M��N�HiU%�$@9#�T��o��.`S��NN�f����,;��tM��>�s��u�ͺ'��I+q��Z;Uï�K���G37=��e�m��AAK��U�[ך�r�����~fw[�e5Ӏ���}Zjվ��&�r�{>S䀭��n�Xg�'R�����^�N%�dԞ��F5H�_4 �q��d�ܒh�8�O�+"
�F(\�;�I�ˉ�ooo�jXt��t{�W�/0	�߲�y$��~����M��)Aj�59 ?j���z~��T
E:��]KtF~W�cR�[& �F����M�9?��K¿$�,j��.3����5�QI4	��ZWݥ�b�$[.aP�pv�J;�D܅�����8At�*����Tޝ��sG������X������9�IB�	����R4F/Lr;��������C�"���ʳ��3<a�r;MG���v#q*pO@K�|�/�+N>>��:nc��y���a__��<I��A�ʆIp�S<�V��Q�7��\	݋<� �^qd.]���x�2/��I��౞���ިq���� �5>z�X���y֍�O���Н�������	�|���n�]����N�@�����www��.��f�{�[�,`8�twU�]��Jf1�����jB�]Ȃ�1���d^m���R9����h�:l����zd�#$��Ɲ"O�/��	�Ï�g���$�۔]˃B�Z,�K�\�ޛ��z=�~�����-����y�G���r�#�᳽f�������V�wI/7c��YQ�rr#�ۯ���s�S��%��~��j�2BK�������*�_���w�w�63���F8f��V��t��8�����P�;���$�R���>@�E�H)M���|���q�v�v@���[����c�G����s/4��-�,1U�����$/X42r>��M�����)�<�����h8_}]��4n	?�&:@'J~�Э�;�eç3;=*�H�wM�]	�tѻ�sB}ͨKK�U|���vh"��2x>^���"^��j�q�c�դU?wӘɎ"O�]��-�Q��=�����ѡ�R=��~��1��ܼV�������:�K��\�%�z+
"����n�:UI˼g�\`n��LTO�Ŭ��e �<�5/YYT�u18���UF\d�>�=�����9g���x���۷�xR�D ��o��n+@,��05B9�U���<\<��gB���o�}�A�b����ݼ֣�No
(�Ե��޼�qM'��镹�>��]�s�TY\�O	&0X��|;�`>!����+z�߼TWɂ���W�Wӱ"j)SE��0o�Ku�!���B}ܧ;!��a�5*��xێ�>"�;�<aO?��v؜��K�[GR�ЛM\C�+O�v�0��b׹B�a�`�4��,ܹ�	��Ҙ�Q�*�;�(�z����(����F�����C.YN-��z�dy8���Ll"��6]վ�d��7�~R����z�:~-��z�ID����c��_�Sy�����S(<~��
 �(��}M�V�K���-���{;A�T�N���f�xGP�k����J�����ͼ�����J��;yR��,�B�;~j�0km4�l����JG���	�y�Ds���k�?�
7�H�u�TI�Г��j��b����(���LQ^��+�F2\9O��l�1S_�c���툎"R��,�����2A�}xv����䝻�O���¨�^dI�4�����|5�F0���U��]d��:����	����0h�=h��eY�_�q_��̄���L��ĺ��	���!�q�ʓ�V����+a�űx�_�)��)�
d��QLN�"YDt��,E�֧�be[���~������3���-Q��/ߊo��D�'$�)f����	t�^�z{}O���wT�=7i�K�>∕��5�b��49�F'�pr�a$J��oEp�Z;u��h?3�kH0��Z X9�G'����)I�8�,��<��]����r��������B����6)��A��G涧�9� '�y(�/i^�S�A��G��u� m,Иm��=�g����a��K�h>g&���8<c�4�,��3�^�CN*)�n)1�3��ټ�� �Э}l���4�[�9v��ֈ�1���=H`,)&��\8��q��|7v�g�{�JK��K����V�4���@�%�g�5C�	~�i1�j��4�.�ok�b��9�0����0��4�#P$?j�9��pF<��l�!���חu���j�z�߷)C[a�d!�1����}3�l��O���r&�<+�c�����d$	��my	0 	z�[昬okk;8?�����r��P�������ء�u���z�3��<vi8�n���H�o?�Q
��>zbG=�L�q<_�v��&q�q��!����9�V<����v�1ת�{}�ԏ;d#�'��3�4�@�6w*d�a�agK���R-�텢����d��g"������O�÷i��Q����
h��^b_<'l�;}W��3��Ry���3:Oc��и�%ڜ���5��HS���n���ۗ�q�S(����k}=���M	�[����sE�F�[#��~�QlD�1��C���Y���[%�o�RĂ�4�Y��+]���=Q���:�:Yh�?��e��[N��(�'5��(��G*V�s,�l���j� ���*.����:�=�j/�>���o��{��:���?�g�3����m��|Bf*TG�Ԥp��}��8F��Q�w�	E���$�d��yP�S�Z�
������_�o��W���k��C��qT��?- **j Y(4+`�Z�D۹��}eJ��9��9k���A�f]O����TQ�勾v��G����B%���g՟Dni�#�d��BX�Km\�3�s����lo�T���v����3����6V4���m~Q%��-.�'���~Y��]�֛�l�Ӓ�S7�xZ���,��d�w!��U[w�����@���->��<���RRs�V&p���zȜ����u�4[>���9*O���R\��(m���ڈ�(j��~�9�ܙ9qy�B���?���9�����U�f.@�a٨���m+�2AAAw��Hk��������*��o+�d���v���ϝ��L��_չ���B�5���z����9xB���xpԷ���LoK��'(鮴NG˰EĻ_2HD�8q1[�"��H��5�\l��@��7I
܋ۍu�{�g��6�ǟ/�顿4:��D#Ժ�x7�&�(WKF��Ğ儞��Z�뼸�����K�#�Tm4�����staT� ryr���Լ"v���9���Q
Ţx���G����-������.<�w!�=��@*zT���k�iE�.����?���������-��@.�Ջ�����t�nP���r;���}�yjm�����z>r@�����_tn[C��O)K��g��6����d*0�V577;,Ynn�c��Z�`�!P�_]�plC[���@N�Sa:�q�)�r��ssy��_���c0�	���|��bx4�02��r�2T�nS���>o��h�_�6����s���ϛ��!�E�t4)��&�G������2��#�Ay�qi�=�����8�JF�n����ֶe�|F�4�"X���	f��n�!�0��_X��
�ڟ��Jʛ��\�g���}���=J+�*���@:�s%̍����Yq�Qi|��A/`Z�8f�N[�<�7���Z��é'yCpp�r��P�dm��'�7ukyB��l���N^���gn��Y4K;!
�Y���rqsA΍<-vW"�'''�����`����dM�ű���ӛmW����K�� ס�� ��EA���˹ž��C�����lhB��~y*���r���zSx���tؔ�v��}� �{{�hw��[怰XV�Jʋ�b�w����?x2�-Yu�!���{I|��~�?
{#�zb ��4{������l9kFYn��h��[DjX��ac[����a�6K���h3^�O2����烠�ȋ]!C����Sd�b�9 ;>������eZ[�3.�w6�\����p?�����^�q�C�������j q�?l�A�u�3������J�ݞġ��Ђz�'����r��5���{�*���U����$T��� !�;Ef'�m.� *0�N��+g,E�S����;6����R,du����to�A��0��w�\��\\��t�[���6ś`rӎ+�U~"�~h
����)�}�->��
pޅ��љ��E���!���n+�Į���<�����m=��q'�$����R�ö%��3�C�i�$����}�p�2�s�O�zy��"s��� N��Ӕd���g �}&�L/����*��"!*����?����p�F9&ggM�W�r.m�re�NjX�fff����; Z�Wx��\p���(/T�H�E~��z��]$���p�n�^?j�
�~��������c�v�;�Y���+tf��kq��}H�!�h��(�H�4��\�����%ǯ�����='����P���o��j �!l�?�tːʹ���	`��vl6���T�������A
��oX9��a&hEma��)L���0M�#wY����C�i�i�e'���ƽ����!W���h�6�E�S8;W���QS?;�n�:��jD-y��/r�76e\��4^^q�(o�R�N���S9%[��vl}<*q��պL[F�y1����@���*����7��oB�:]�G��) ����3�x1 ���Q�znz0�Ie�^%���J�(�ງ&�M���ْ;q�^K�w�ζ�+V˃N�a�-Q��w�2b���N	��L�d!��ąnɉ�hҡ���bd.�e���ƥ](�~�n�E���H�fiV-��tT�u��ψ"C/1�齊�]����,8T�۞#�ፎ���=����r���(>�B�{4���ͩ;Ù>ِ)�)x�!�P�B;<x�=����^�A��BT������àm@*0ğ/b'":����Z��g���Й�Q��hr�P_�E���y�B�N"8�:�%r_W����|܆���Ї�!W��BF��.�����Q��Of���|h&w�m5C��p&w�_�p���#�2~���:��O`�Ԍ���r���K�Ha�ז�N W��4b�d��-����b)o�E"sV[0<��'gz�8[i�_2ljU���C7t��~��|���i�/��a���p5������Fi�� nj59ԠE��#?c��J#�6N�6�Rƒ�'s�o��X01��t\H`d���"�ٿ��Uf�kl�!BX�����ܿ�S��UA�V���^�MWW�9P�%���B˵`�_n���tO�Ӷ��:�_����|�j�01����#s9�6~oo�2>c:I`�o� �ɄH�|61
��߅	��4�y�����\�C������-��k���ٶ�L���}��6[�M�z&Z/_���%t�2P�LP��b�/k�b�9�Ţ�^��F���i�v�0�XC�~f.]���m�Rh�$��8���uϘ�z8T>�k}ﻄ#Q��$�w�4�TF��ǌԽmy�v�R� ���\�:�acccm����0L������鸑zd��۶Q�fG ��4�"�i���{�@�n_LlJ8�2R�&CS��"u��Ö��t�X+��
��� 
Z�����,��v��r���NJM����1��&�0X�n"pђ�����|��*�+f����_&�m�L-�?�e�}Myq:-���-Ow��}ኵ�Q���IkSG[8�`���Q�i���F2��l�8Up����r[�(��Q�Ǒ�w��v+��iI��B�o8��0�?�� ������I)��[�V���d�abSp��
T�I�}Ӄ�F0�c*%c����Ҹ�˅��;	/3I ��=�D7\�A��?'�/��mK����me���&e"�7ʉ��h� e��r2��v^�$�0'Gf�2 p�6�,��ez�P���1I
��i�1g��:kA�<K |�W� �F�D�6�J�@����9�����=�N���������z&h�Y�����Q�����n�[8�~96�~Z�`$@�qy����>��h�ݪ4���
�Z�{2��W�!Ui��|xl%~JY�g��}4$�~h�M�s�%��@��L�*A8���8�^φ�d��
�����J�����
M�$�$ ���YR|���N{G��`��-Q���`Z��o��kSO�EN���z��`错�%����RH3
�����H'�2�L\���TSC<��'!�/�QĠHקa�oEd?�>=y�����佝��2�J�`3�bS�T:rTDh��	Q0���i���<ĩeտ��a��;%!B�!A�WYL���?��e�8���}���P���Gdѳ�m������4��{����E�����U�~BP�f�5G��用L��G�3������u�SY���Ͷ��˹u���$�v��6�Q�`i�0���]�U���2�hr5(�b�"Z�^��]H
qI�\V�����ûu����J$
�������H��ƞ�x@ҕ��/N
�a0gu�RӼ��7�20ۥ�j��O�v�U#Q���ۇM��u��̴�5�5t̝b��𘜙�|�>æMt&y�Bh�;�x*�r���D�Uh�YEM^�i
r��\�]\T�V��S(�şt���<�T��8�IU�,V���@1.�{q�7n�[����(`�އjq_ �^U�J(�h+�wu��ۏ���7��J�F�.�%��VZ�EMS\�Jd3���W��7����9YI�'I3��"I�,�C�$��z"�&��SsB�nߣx��IW�K5�M�GT�nmʯ҉��Ө%�C�9����,)l��!3�:�՜*X��?�U3��À�qIJ;n�?\�Ux�I�|cm���ϛ<
6�,2a���G���������a��h鋡������Y��G�`O��.��@�}��x�|���$Y�GlniAI% �s�/hH�R�#�j�sȴE����!��tLF^���IU���.���={h����+���%��Ă�HX���7P��-�YRkB�f"���w�c�¢�\�V��
F ��BIw��d @Fi̥��6�;=�Q���ɏ̒C[� $N��YK~�h���vbp�k�����ץg��2�V��a��U��&���U�k��+��v��Pv�l(����S�P����<��Ce��6���z���"W��͋�}#�B�ъ��a�+����F�Y,�Tt�ܩ�yr��
��W7 �m�gM+�}Lx�0�H
x�<���+���y&�gz~�2��Տ��C@	��O�����C������K')E;<���M���_vZ��MxU��S��u�p_U�n����M�M��2l,��9c�P��j3�|�":W��(z�;!���,s
��ٺ�:�M�]�,��32Xϗ�⭟XNd���Vx�i�e�[�8{�*���;4+�]�ŕ]������4#3P*���t�{�zs�q��Cnw�$f6����}���W������\�r���GS%�ixEqȢX��Ey��,����!Ry� �`�#%J�����cŢ/�J8�����9e���F"��G�谘z���Fc� r�����x����
�s����gXj\ઉ��r���>1���ܩ���S�@��E�ف��o�~����f�d D)��l�5+��۾ �ߦ:���nnn62�ֺ��/��񢀉��-���|�.���`�㹲�f�c�㲆ow'��gna>�׀���0
{�An5iW�����Y�ɏ'�:{pb�����������N�{�n8��#j���2�&��-9�0MLJ%��I~`��:W��(�/ ��e�TUgKu�-`Ђ��@��V���1k�k]Ɂ6�.\��Q��DC>@p��߿�節��tnu���Ȓ~-Iֻ2�G��u���g&u���RV���C�ͥgLi��h�F[�:� �%�ʪ���2��'��eaF�l��~]�����ϯ�b�nn��(��n�	�'<Y���P3�H&�0�!a�,�zҎ����!��_�wϢ���o�9hH)+&ѥ�
"0���OA��^�?!�w���F�5��|�͑jo��DT��q8��p;5�����M!�r �I|���z�� l֜"�������.[6����~��sop���С�~:�=��	𐖖J5��顈��	�D�wL�Kkiiu�8����>4?���l�!���-��s2�"
��ݩP9�/�!nA�j��a����ڔ���ͯ�#,�!�0�Bg���8�����aS��\ %�~NY����CJϋI|(�B���׍�Q~t1X�M�-��p��5�֯1Ɲ�z�͞�&�����RXd��:�A�Y�-B��̺ף�nޟ������ED����G�u~�(ذ���}��DCC�Bk<d��%��l��%�����Ν3y�W��� ��tf>{��,ʦj�D_��L���4}����-��S� ,i�P�K�PL�$�?v�J9� ����ƢM�Od�F4��DلI�=kOH6�R�E�DaM�Y��GT�c����S.����m%�Z�#,��N9���z�B��%�ہ�՞�'ˈU��T��TU�?�U���bQ�T@u�Ä8�EIL�+�w,d�R�5�7/����2�����	in܎�'NJ�噠}���:I����k�����.���*��~��~´"�WjV�שj��XX_;
{/��o>K���Z����%RA*�ۂ��׫z�g���u]Y�0�NǇ]������_ -�a��l��9|Gq���Ɋ��D�����
'�w���� 	�>#:Q�3`�CP�I��;a$j����ŷH�9?W;EZ��D�aE�*��*�n�������q�[��W��=Y/��~)q����P���x{�ӱ�2�U�D�o5�x~�ߎJ*�d�G4�J�	iizWx�W*B;Vh��FΥ��ql�t �������}�;-����H��9Li���p\�d��<�|#���֚f��X�]��b65���h1 m+e�1F�ё�м)� ��p������IKe����;S!b�Ǽ�P*\'��Q�2�H!�y��u�\�ßrt�
ᗚ���I��܉�m�^N��*�r�>/�>*�b��"o��� (l��h7T��!z��*z�/��T�����,"t�r��������>'�sCY�F�"�az���o��lF���}��+�+2��>?"p��M5bN�L/����'��ZA|��f ������!���q����͝1u�bUI&:599$]Y��|~��_�^?�_hgM(�G�ꦊ��q���d�s����'����χ!k1)��S��?s��?1���#��϶�%si��w������C��x��Mt�3�W�}���S���z���)T���蘪r����p=��N{��(�v�w:T�	�T���#�
qi�[|�����t7����W�s���0|%�oLD�AN�����\v�<�]�a�)������Nu���+`�oB��45�C��oڀB��/C�w�Tም@)b1 ��
����⧝�Z�hL�Ħ��)nJ�%�_�r[,1U%�2�T9T�cgU�	��jJ��|�ā�qJ
�s�T�"�&�	'jX#0�z���F���$�^u��"����,�=R=�g/B�����0��0 �e�*Qߋ>Þ��I�U�2�k8L�k�fstiD��}x�%U��rb9��𹗆V�@�8 `����ІV�1-�̈��<>=9��j1����@kj"��__��ȴ�\L�$b�F�c����k����no�r�P���6���$�?��|\1O�:��'���8_���,'�
j0$]�3F|D�""��BR.�7��lܛ#p��)$G�.NR3}����ӳ!y��<羠,9���_4〟&��g(J���!�oU'I�"G>���~CP��N�1EhJ4 �I~?+^u��X�r������N��Ir@p
"�K~����C�pT������������Rs��d��Q���%��Y+�zz��g:�zV����R���_\�	�ˍ�a[a����SQ��y_^@� �2G� O��:qv��f|8�<D����+x#�o�t���:(�<��.`D��k��y�[����S�P���˾�u�h`)���Fm����L���2nd��;SK������q�ԗ�d��a �`u/��/V���/u���oY��l�Buq�}�>QӉ:�K�R��-�9���(5`����'�cDK��Gt]	R� "xR�a�]F&i��T'���g�PY3X*Gm�f:��~� _ۧƝ�j�u�|��6��{�K��:=;߸~p8�	�6�+kao///���PB�]
��dBbf���P<��2�	��������;�z91w�o<�gq_j���(�C�0��?��,rB#��h�s|x6��Fɒ�֘�Q�S�M.h�L�°eW���8ex2���9�~�a*u��1��37#I%s�H�c;��|��O�1d�z�������y]Av�ļA[XQ�����F$���}E5,m����d�����XΜb�]S;��̶�5;�2��x�3���B��Z��V�z�~�sւ:��3�(v n8�k:v�u�B�������y]����]|hZ�K��%S����T���~h�f��.��&�v�@쏎B8C�>�H�j����O�c����ԓju<~y�"���x����~���%���y����-�M�ז���#��
�aCE���NE�MU�hHNI�a� R�ܐ�<Wi����I� �S�t��8��>8��*�rfk��<��%j�4��45���$�+)��T�9G_i���H�ؑzP%��DMI�0��a�����-��KӵQiE�_u&U	Uk��T�.O0L�6��iL	y�i�H�V���W}�>���R��~E�w��V�� n/m�z��WkB��N�Q����E\��I[t��ٿ�N�07�?���v����)���e�+�0X���gR7���ei&���Ɲal��&۵f�O���{�pw~���y��4~�D��	���������y>>>�ۣ�����Rg����zT[o2�ͼ��q�4�y��N��x��eFp�\���3D��5�5�t��:ͯ�|��K�lu�����^�7'��=W�Eu�-ӹ�~ϨI�n��2U��}'h�t�d	F�om|���+A�i�D��{&s��)\�ў�a#SQ�9N+�q#�k�W��H�N��2sQ�=W���B"���G
���.�C;W�,^��K<.I��ē�bK_Qǣ�6W�M[}�D^�S�MԪ�h�蚉W�U�}�t����)���I-�npCh)e��s���	㆞:_�ܠ���5{�(�{���ф���:�q2���<l�����m��G����y���qa���2�
�Ӌv�>����9t�
��rU؊;aY��:���w���2t6���P-�7�pf:f��L�sro>�������[o�e	�uz��M#.�d��!���|�I:�y�ꙁ���2�I�D�i��@;i��%f=`�t��@�}Wq��?����*yc������+��pX�Ӿ�h-�_��#`#�n��!��L�G4��u�A)X����&�J�O�MƸ���?\4O�ٙC�jOb�C-����Wf+�I���U\��F�u=4RBZ�*Ն��������{�(�_�x�Xh*��@P�Z@��8�տTg���q���J��[$$=g��s�il����ы�]D�H"Vص���)(�p�r��g&^�$4r:�C�g�R�SWI����L���a�]�8F?�Ixc�l��5uY��vtF�w�;b�
R��ɓ�h�ҋT�?j�7%|�1�/�G��ni��L��'߹�N_H·l�I$�O���aZ�ݧ@y�,_����˗��N���O�~�����/_$ͯ�=�-g_���U)yn�0��#b�@�j$~STTTh�S
_�vk���7%]6t�U.䡥�E�S]�?��ww����D��f'uہU��f�5�˅��a�b�����)g��nV�P��5����E��1�D
����xQ�G�LM�G�x>l��"d8ZQJc���R*�/�;���T�K�s�`��~)�e[�4G;�H��h�F�̘�sP�q����Ôz�VB���,@i��Ό�(������P�T�˺|o��oh0��MZ��
^��/M��5=��C���q��w���vI0���ri6�k�H���<\16��V�|:е=p�&lٟ.״H^o\N�^��x0�����1��Ù���ޗ�B^X��k� ^I�n��/[
�pD*�F���߱�4j1"���Wɔ ��U�1���
���Ɣgĕ�C$-�BC����� �5d�d$u��@ 4��B�:���\�G�-%j���]��ci�p1�R�qу1 m[�SC_џQ*���� ��^Fm/��v��!��*���rj;i� �S�ln��޾�Te�����nˡ�g�a���?{��3��P��pPBq�ɯ��	��AXF�z4r'Xc�]�3Zg��$�r=���a5���M���z�$ܗ�D�
�t��A/�:�
����ycM*����v�x��i���z8}�O�%C�׫�liZb���/��N8���K������`� ����o�ֵ���/{ci�:���\��5�u�8�n���g�����?]�C6�Z�w����&�*M>�D
���=�L���a��`(��M#Tc�����E�[Vr� )�@�"YE|S�`w��v\�]��ޠ9w��%X�M�I�9�Β�ςm_��{������s��.7M�*m������ۄb�1�v�@�T�����b���V��	f�����z��'�T�w�q�L@���pY����B��4sRy��IypgZ�s��i�w�&(&���霵����ÿ@�9	#��=	�p�q�̀�H�K��j��B{�������1ּ�Gy�)��g�p���2Oݷ�L3�J�������5�'[(2� �ğb��[@gW׽�.?�I��ק�z�ezc�R�ں:��LI/;���	nD��j����j�����~%�ؓ��Ģ�"Q��Uѯ��^��.T�l:46���!9oF������l[���#��Ǉh��~Q��z��T���A�_.�S��Z)*�w�q7~��1���I������iȧ2��zu~��ѯ)RˡvgO����?��rC.da>���KP#E���.h9-���d��_L��ɜW �U����z*¹t������:�������\SZ���(0/��!x<�������;��#O.���%�����5�Kݏ0C�PW��y�qx;J`q��a�������V�b�nզ����tb�Y{�9aO�V�����	��4��ja�J�^<��U�E�?}��4���EaɖЉ�O�[]��e,L���;IsN9>�l���]��׬X�,g�p���D����df_�A3H+:���$�{.9���a����W���>���.�K	��嬹�\�#B���8��r��P��$�����H�G���O�d%�P%D����-�N�U������_�K��
�_,��\;���д�~�۷�LQ�d"P)>�$ KNk{������.�����T-
x��������0xC�-Wo�:8O\F� W/��'T� FQ�H�:�viO��XXO@�Md��`��Da��`�Ŕd?�׉q��E�&����.9�q���3�����-�ѧ�Dj��C�j�@���1sq�_ox�E��s-���ѫ�yCp��O�7ύ�9[i�v�Pg�������!{���,Й�JLć�<�̕O��kЁ,��I_�l�㱽;(�XnA�~T�|�.��S���̴�^��?'�Lj�F��Fv����ʿ4C��vZp+é7��{�YKG��:YKP���h��%8A}�������sp^C����ƭ���Ḯ�c:�F�� �1��y ;A���2��hӼ*��*�Wb�WV���<���+� �x82<D@�Ld±�(���j!�<�Ӗt�d0j����8�B]rְ1�A���&��n"�N�q�DM.O`�v8�4z-�
�5P��B�+o�7�:5��I���.q���S*��aZ߬��K��q��:D~^����о�YY<�GN��̻�P�[��j���ލ�_H�ځ��*^�1Ĳ�w�kelw��������ߺ��H1�j�X�<ϸz���p�2���Q�EuN4-�<���ܧ'��{�%^�>��'���z/]�'mnV�������g3SS�8~n�@�	�ޗ䤤����v��Z��;+��tT�������ҒpR�]��bē17{"G�ӥ����U,��p/8���F�jR��,vN7�`xr+��FRW3BƱE��	O)���I��F@���,�ŕz��h������)�n��G��{�t��dc�i�ݷc)��@_�]�k�N�B�i)�T��o0�T�����e��?/|n;��c��J�C�r��*�8��A�y��S��O1V�f\���c(ݶXgM�n;�L�.Wlal��1��ri��Z�^L{
�"�E��ʓ��l�,����]fQ}�Sj��׎n!��K���~3����g�Z�_8g�8��m,�?�kbYXSf"������/èE��s�b����p�/i���Z�Q��Exnb	3#~*����}Ԣ(Qr^��W\}U���;`m݀>a���<���(!��K�H�yN�����u��^���R�Ux�8�P��8��n����Ob0����Q�~m����v4A~1ǭvS��υg(Q:�I�;'�d1����K��h����f�p)�=x��s��,3Z�l��Dѯ:��:��
����1xv�ĺ���Sㆇc�?zG�7�� ��"U��9�qn��X�O��F�*I\���آ�+S�Q�F5%���:>ъP�<�8".��Œ�(��JЫ�Z�%��i���gg�O(�k�8@�x~0�G�[�KZdD�7"��>���~�o᳡sss����\&D�Ű"��Z�G�A_�*�ڑכ���[wu2f�:��j�m{S�q4�{�Y�vXyb��Q4q��_��'}\1$4����O�d���$6���XA�^G&D<��D�r�\��S0d߀� XT����YDS�����;t�)��	������m��������Qv�V̂#C�e�Uw�_
le��Sr��"̨��Iߐڸ ����a� _t#JJ�97>���%B&í��tN��+�YC���TQ_�'���:X;F��ֽ|n�1j��Ϝ��Դ��ȴ�lg=a��Ȝ����~�m=�Ȳ�mN��9[i�<$����o��l��GB�vo�\"�b�j�T��Fߘ���FaP�Z�a�X�Ec�;6,m���M'��G�䚦EA6)��-!����&������@�%$}��xd\w�|z�v��aEy;,c�a�Zk����9��'��XTqg^TL��U�^�����R�� <��W�%��9�B͆R՟���Ҕҍ(�_r���<'�` �h�Np�7��4������E�d��*���2����z��8ǘw�����U�y4��[g"ޞ�uӼ�P�߿I�{��qF�+{�J�8vzۺ���o̻嶘�s�HʷP ����o�����òb>L
�L�e�~���Z<��-8�K�ڐ�Oѽ�l!�'(�2K�������Ѓ�g,�QK�j��'F��,)l<�0���1��=����5��CnX,���?��
��DP��������i���Mx%_B���`�����
r)w��'�}9%������-�B&����=�h�;�L�"���.ZJ,;�VQ����M?c,[l]\k)1/�q���'L��F跸� �[N��a�9R��R*��r[ZZ��u���"��z_,UnI�ѓ9%u�M�%d'D�#�3����{L�>���	9ѯ�o����&
	4�F*����c�
�i�B���/�Uq��A�!3�1�~�NH�\a*Z��7z``"֊V� c�`���
��MG�9|���-���`X�wV���m��ӟTEm�|\���	������Lu��Q�Yr��Иց-�ɨ��8ˋa�;�Q�W��,p`�w!G`��(o�+��uɴ`��9d�V֭�
�m'+�q2�������Q/�갋���\&<$(W1��~��
�{E���K鸦ͳ� ���[04�����(&t���Z�r([Yl�]��~�J-Ϫq�$�Ԅ��\9/6B�Ụ�]�>������vY�3�{��1a�m�q 4~�2 �A����d"���)�'5JJ���
��͜���앣T�� ��ɻV�恙a�� �i8}$��!p�j�UF�⻼2�:ϙ�o�Tp�ma� �a�;�@mN���܆QB6�n6�E ��E���Z��pL�5\��c���:O֠趔��V@�k{`�d�Bx�a�Y�jdk8+8qo�v<�K�����B����,��N���w�AA������I��0]7&�������	��C)��2-�{#~����{�ap�\6������1��(�܄%T�R��{Ј��,e�˴�x�d�`}��B����;Ǯњ?�C�O�wU��kBX]$�W�1��{���T+��d�Ř�jVlg�V�u������)�`̟t~#�Ɂ���*�l	Y���Yp�p�Q�0? �����	��^0�C,~��<P�����&��_x���UU|r���smy<S��io4��Dퟨ�Ɵ��А>
��ikk[�\��E���PG��/A(�����,屍�6bG���U�P�^Ma��0��S*)�	��Ԍ��?e��RCxrɕ ����Zb�"�}�*�A�W<<e��s�?i27S:��!u|�x4J5�G�A��r>	�3�BRX���m�)0\v�X�Z��qB����s��l��`˩+JZ�q$8��q��x�+	����4S�e¸a�uܺ�����@_k�n���:�I�R_����0��CNnll���4�7�UB�T�w����������/��:E���;ޣ%h�,��"Ü�j$�K,��}�S5)jt,��Ag�:a?^�"�D$DCЊ�4]P[]���N�X����JqwwNp+������݋[��.E���7�3<�a���{�컻g��1}�ЈBX�܎Lt�+goK�E㣋��:�4�2���0)&�ޱ8_������ ��3��zG`OJj��S���3~��T��dA�)�d#��%�7�mX�Ǐi��' ���,H���5��Y;�[�W���t�|�O���:���E>�_%U�o�<�#�N�ܞw�k�Xf�iAQD�I�Vz�g����Y��pz��~�i��w�9�d�؄m� {R)�Ze��3�s&��|����Q�Z�抸\����
�]#v��#M��<Q����.��;οaO�A rv�<��a��At_Gh���i������V0�����vHx"�o�swU=B�w�c��&������yƟ��/�!+=nO�M���a�S�����J��	��o���J�+<C4�soi�y�.zCCCO��U�R�/����Recә�-����?��;;�U�~�+H���,c���c�(��U���i�y�,�[
�Zh���W(�gƢʠY{�#Iʧ��;�3�Y���.�����~0:j���d�E㍺�rq�X���s�(��z��%L>��)H*�C#iz��!�q����})ؕ������x|�����v`���H������@Q��mr��体i.�^,,F�����c	��յnW;��E�2�ʒejK/�(9���s�V+E@X[� �����J���l%o,E�=#���_N���}�U��Z	~rB9-�}��tB��W���SV�axTtpQa�[�v�;*�Dݑ�c����'1�5sT���Ӛ���$.�y�y��L��?�xxxT<]t�RRRjԛ�1��0����P/;�P�ز��77m��teΛ����ل�\�����z�z?���p��J�~��Y�y��x���4����媗>�؋�U,vv��|y��G�w$
����%ilP܋��;��c2q�3�~'*J��2��Q�%طq�4���Y`�� �0�5-L��s ��Z�Y� �T����u��ʟ����x@B�y)j�G}S�pߏoLP�8���O���mن�@떡�=�tN�C�,�þ�f��\.lRVXԲ�
�z��O��vc{Rt��5P�N8f��� o�>!�������P>M��:���M|h�����P�IH8ڢ�ȉѧ���;NeD�U:�P;.\m�,Y�a)�Eˬ�U9�
�a"5�E�bD�B������M�q����~I��d܇�����Z�[@�7f�Y��[H<�ص����O	zD�t�L���6������g5�)�ݒyt�����[�l�	:������Tu����Ǚ���k����ϣ�3�f.m���r"*�>]fE�7�d*o%�Yx��c�Cb�����(�D�U�8��X�!���l��!���Np��{ؕ?��0��N�]˘(�Q��ڜjo"��.b,�
����2/e���'^�ځ6�>]|��F�ʩOy�㺜�O�mv��%p�.nD�s�eh���G���8Mr��W�4�@���:>��'
�g"s>�G��㤿���g:;�X���v=T��RyVso"������++�ǾųN�,,q9&��s���_*?��QIߎ���tlg��������5֟WG%׌����Z��h�=�f�6����k�g���/����\�Z����[�4R6��Vm\��y���uܓbԨ���1���,&�ڊ������;)!��+�ظr�o�l�*c�)ރ�NS��3��'=�_�(�����I�q��u����2P�|"��1E{�@���FOwg�����|/	�5�>ڛkBw�ꗿ/^��E��7�b�7���?��:�B�����R������3|i��VJY^Br8�w�C�ۢj�i+%��_"F�����cc�+{*�9[xf"��JR�¯晘�?�ޙ��!��)�'�}�� l�:+;���q�����c'��%���5)禜��6���Sl}e%�2���L��H|vRP�g�@Lh��Y�̀���Wو�6�u�a���;z�lhS��uu���^�(�(6�-X~k��D��1^���#7��UaS���O�+���������T>B;��5>k)�Io}��]�bC��#�$7ps�^�\�;�k-+C&��?T��2�`����Ӝۊh�����t�om�9��:&���F�o	c2����)L[Ƥ$�E~m	u�*��'���)Ym���(��T����6�?ړ�ՑB+ۜ-w&m9.{5j��_Fv��w#��O�&,�Փ0��#���]�n�#@{z��b��\�lkû�/��H�,��o�C��BTupå%��NF�G4���)%��Y��`��Ji�
^���Z��	�	��#6�����6E`[�d��P"���9-��_��%2���0,Կ݄��^Ƚ�f����X����k�6�~�lj�,���ٯ�4P̵�=GC{\�6��J3�x߷��;��ݗ��e�.4�������D�lI�5�1�����=&��h<�]��IF��YDCaq�st�?���a�k2Y�Z�������멫�O�y�a�����>����>�u�Q����G���.Vj����~N�'���F�6=��!����ULD��������Z�\���R�j���=��ЮҶ�Ʉ�L�>�����<D��޾|�Õ�c�Z)ܚ�7��G��ŀ����r�fӬw���5�И�]����� Zl���>��݁���������y��1Ru
G�_�01L����k��1Np��W\"τ��a�T?ey\Q�ӕz�Ơ9��'Mge0yM����D��0�<�_{M��@f��V�vh*�	�Q#��'F�.bHtd~�k���$ä�ץz����rqj�;1��7D<����ߨ�,bd����'#��J�o,�m{4�d
g}�_I�H`���/�my�[s8*L�o|9�hw�������mG@��� 3N,����(�y�Q)�כ�v4c�g��%}��F� �S��ĥ㾗xxr�o���N��7s�|�p��#�#��-zh;��g|hub���¢bV�͎8����9ih�#���qX���|�Ǻ	�$�����P�ǽ��� !܎-]!����u���{�!�Oc�3nwن�ҷ���MN���������~0���t7�X������m�eґS��o��=̹�������G���%�Z�QV��u���2�w7\�L;d^��x?/g�Z�?.Vh����;h�K�L
 ތ��)�X�h�.d!(�U�7����e����V�K�=Le��	�݁��C?�І�VԼ��������>ww�[N�q`>�\k�zm0ⓓ�"��A�����~cq�L����#Q�k��L1G�bB].�r��B�j�e
������ tX/=�>\�ԙHn�{$�m�2D��Xj�X}��{ڟL�:�����uu�7�cZ�::?"0���b�m{�ɔ��F7��n����Ѹ��Y�ƦEX���f)���(s���6��y�,�j��h��[M������i
ѪI�����D
POf�i$+��E��$B���e�C�}���z�\��h������}����E�D{ME�Q.D������~M���4)>�g����B2b������ {�;e�#�d�\j���九�zՇ¬�Yk�=w���g
P��o�m�����T������-L� ����,#Cn<l�� �]Ո���-7�=�[�~]���x��R�@rx�Q?"�����/�m��T�^'�Ќ�E�5.O�&b�eX��W�;:ΰEpm���S��[>C�]�3�P�{�u�rO8��9� pY?v��\��],D;�Փ� TR���E��������r=r�\����J� .o[O��=��Q�zQ_O�vs�\�)�ﭳ��c��fc��ts�Ծ�ab�2�h����r��U�����q�ԃ��_zt~8s�+��vRUn��3\�n�-崡�bF�\mj\#0F/��N��N�-W��AOg>�먬�r��Κ������0�V���9$ٵ8��¨��I4�b�lDN�;�s2��E�'��������~�o�h���*������4����9����ׄ�}�G�	���薕+9�=�BƔ"��Ⱦi�E[Y�mˠ|	�)KI�V�#j��1�e�Q�;s���`���@.�A!���:�M�7��˳�*���������]5����O�*x'�f��f���-^�����yff��A�k�@T��̌�]��
�������FG�>�o�F�-��^�����Jn޾�� �pf��I���NE��{I�?�c�c䜮b�0��p� h��Ą��  ��x��n����C;"��ߵv)@�蚥 ��#�M���OF������ ��/� �6���?��\2����p�v6��&\Q�s�3b8���3S�O��-/́�c�*�	��j��������9>3Z�K�M�u���~�7�	j�ŝd)1���� X�ЩJ훓��j�[�fޫ��K��x �k��E^t3�F���C-�^��L��q��	�'<�=�|zM�"�%W#�1	.6C�~&0W��"�V���aO�\x,���½��	�,L�I�E��Ӻ)>��1��%q,Dx�Q�w՟@<w,�|G�Z��l)�0Z��Q�%��gX?��X<Y�3r�
8�H80� Vʙ9�1N�Uc�U�4�H���Z���r�j�G������$�9��YW�a�l�ӂfs�>�\-��\���-8�A�.P�����ؼqد����������)2Dj�B�$5R�޹���v\I44�Q�TCg-_�jt�x���e@��������� vNti�f�G��5&p�d�C�dl+1�zUB�����=�@��O�����T��Gqx\�:����� ��+j�;�v�Z��o�X7��3?|Zϖ�T��ph���<�p��p�Pn��G�>��(�h��,��J!�͒�3��{oB��sJ�_��}���l4g�Ξ�!='86.jx\�� ���zM8���������D����Q���a� V	���gXB��M�Ĥ�uZce 4�?����1��bJHH��r�}���u����4��X�7G�n>�Y.�(��[D���M�������yI�~��P��ZW��0���Ѽ���<B��Ub�W��$���yj�ĕb@�C�	Ë�NB��}�~�-�u�;�C�rc�v`$j}M� �l�q}�ςI ��kw��
��B�u�@�!�K��{�]�K,��4D�#s�N�:#h�JlU���'�- �>�Vi�=R�n��~����GBlw�9�{�~z�1����4�Qz+Zkd�����bZ����ԭ�­4�x64�7ƺⶥY��/�!�Sճ:2�6/b��zډ���O����)T��w[4����%� ��!��~��}(�zr�S���B�$k�z�Ju@x2V���â�7@�Ӵ�'���yxx���Ճ��^86=/:�&k�!�3���-������kn����0BI��N��/��̮�5��K����̚d�#ʁG�%��^lP��︯��۬ث��~�q�˚�Y����O�[����l�p�:��������_QY���ļ�1��(���]�B�Z�%�i��o��@��~e?%3�ј�]xVb[�o\`ڡ�/�}��ήC�{�!Ϝ�ZڱT����Q?5u�3(l�]ɸ���=��[
�bO�M�û<�n�#��|w]�a#���D�%�5'A�kv����'5ޤŖ΀d�G����X�&j8����6S+a�?K�:��;��0s�^.jM5s#�C��{�_T;Ji*�m�4+��Kc����z�Lrw@rF�Ȳ����IY���N�����r[&�?u4�&>6����Nx��0�ɭ�O�$&��e�m�(�BϚ*�h��V��=ծ�
rI��K��2��������Z �X�O-~}7&:c��7�@����CPF�X���lI��H��2�(��ð]�?f�@��yVik_���71�<��Eë";���߶c�@	�E�$��uk��T.��߲�Y��ӂ�6����[�\� ?����}4nt}XQ�*�pIF�u�X*Φ4�q���ډX�㞿.ZCT`��:W�*>�vUO���뚈�Z_��3��mOJ����a�Dw�î��t֤�A�0t���C�r���sK�qa�1�Q���{���o��й]�`�(�tv�9*��]KC �_40bl �1�߾ZqH9���u)��{�����3f[/?����1h��Ǿ���Gq5��������*�lT����4���F��yD�(���<��S.q��O������\8f;��O>���U%m���BH�*&:)�%]�lH���Wi��vȰAPX-c/
۞�`�T���B�A?�V�ә����|i �Z,AG�X�88�B�bH}��iv�}Qn�Ҭ����"�K��s�v��5�'E����R#�Ƶ���Vy� �*+i����̓w�p\Z���x@cr:/���@AM%Y0wQ py���I���G��m�S���o�ڂ���k+b���1�S�A�����9P�A�/�������a���B�ŧ,�)�iJ��SR����`u23'�2I3v����,v.��Wy=�8F5�ص��	ۢ�y��(���>$f�ASIЂuҪWX��л \������bM��akR���m���n�A�Q�D�j��ueMj�MKt �j]\�Y��;�Nrt]�6�տ�{��HO@/�\��_��o�����nO/��@ �M�@=h2o�\��M5b	��B���ͫ�����o9�{U��2܅dU�Y�RƲ�Ñg���$�Y� �����5�_�.�� �Y3��7<��%�8)׋��U�Nb��ʭ�Z�Gp	M�_��s��~**Ρ^���LOM�4�����Hu�a:is�KDq9���=>��8)�ݬ6��
)��6I,0�q8u:�8�� ��G��x�R��BW�=�� �1���i�36�cX&�Rh[���͈��`Dk�� �&b#�+��D��Da�l2F��(Q��ȇ�]g�V%����o{1a��}��C�}1�<VwP�2/����d�35�+V��~����P#T�����9a�m�&��t�� �F���IAP���8�맚+đ�|�'�W�w��{�^7���wi��N�I�aV�1�BD�j�3��E�N�q���-]�BIT�Q����jd��- �o
�>����wM��dce�4�\8Z���96A�1�78�̹��ᨊnC�Y,'C�&���w�`+l{}L�P����S��x�B��ڵi�K15�^3M�&`�9��^�0蓬3h`q@;����g���>�"\B��o�ܹ�}����Ȁ[���'���۝��+��ur���*�����[PG�	����7�L����-`���� ��CR���7)K�v׋��t��ק����h)KFQ�X���T�L>���>݆��\��qQ'�U,^��^��*�I��[xx�!A�茬���F�(�����(�����'�O�|j��Q�����T���yv�௡�����CqY�y�q�7BJ؉S��������މe�-��1�~����fRQ��O ��C��s^�L�W�U_�q"�s4��0��%���2x��7�i+��F-� };s{�|#���(=8~��$�����.��.~��1����bw Tq���x�C��"�,���z��5�'QLT�֓�v�,����$�Z�F�dםi����Ƙ�P�#�VQQ8M�����"��%�5�@����z,�):	��'HrP+r������w�mpK�r*Ms"#��
VSF�ێQ��/�#&�6-�~ѡ��?��;��g��~���l)�w�	i�}Fv�K�A ���۸��d*�c�IH�w��'���t�w��M�CM�D�;��>��>��:��!3�!��Q���c2L5'RX A��/��G/T�(F�m���("�A���Ҿ_f$��ƓiL�ņ�*a��1����O0��0$$�OT��_f�I�؉�ᓪC�j�7zbWp��6Bql2���tZ�Z�8��vG�N8��kR���#&�MN�I��R�c0�`#b�}����	DIY�QE6)���G�JH-���:R�!`�%1�=��ի��a��<���s4�l[Λ��M�ǃE�o��S?����˯h���`��f9��BKK۳]���GP7�����.��!��.�QeUU�]O续Y���M:��i�=0�ĩ�1$LH��bJ�%�6mN�υL[9X�d܊{3�%U �^)�o�ff��s�E�Jr$�Qr�y&!H2�9���r#�:6<�Ut'J!GǨS-4k�{��e��� ��>Y[&�C��غ>��D�����s2��S��?���k�����{����2�t{6\aU�6 T��f������|���\H�	�������˰ƍ�%�����ڼ���ͼF�,|�|�2�YlX;dPv�ǽ䎻U�R�|���A��؉^e�f�"K��?��\�r�71[���JJ�5��kS���2)ˉ4�v3�M�m�Қ~�=~W:8Y��W:�u�YE��G�A��<ġ�?�z:4Vm�5�a�7��>�(6�D053�h�?���>|f��� l"��!I���g!!���tdI�W���Wu��z�-$�Rnv��o�� �ɹ$�_}�<��9�Kg��'1��6#�wK� ��#g���/_���pkxg��
�w�/�~�{_mu�@I��D�;�̦2�@�U9����?>��T�+�C�Fq�]���D�r�zgog�����A����[���?V��k3���w�MX4~]�M�%�o�>�	N��f�<���!fQ;���M�o��)����Y��`���6vO㧈ڀ��o�=ή���}�.%G ��(U��6�6m�K� �:t�5Ej�k��Ҽ"��ނv��b��ro��Ǜy��s.>�j�j5t�o�'RX�?���7#��H���Ug���r�Ў��:�R�咮�0�j~- �g��=f�ܖ��u���i��0���B鲯X��[��e_1A2�$����I����r����T+++n�$��9e�w �$SEUՠ����о>QF�k��P,J�, �ʊ��(��=Q���kPo�m1�7��N�x�0^���q�iܷ^��}o�+�Jxt�)��)��</^#�E�C���-�
��j��͵�,�O<l5_��G��
A2�4	����6��&&�	�
�̏�#�)rZk�U�Ց@&�'���-k�00��u6	�'~H;�ba?��;��������RІcE��J����eNQLɶx��o.���zۤҤ�үJ�_s7�CQ|*��z"�r��8�E1��ZcH x��	=��ꎗ�����PP�O�� ���-��]|�{%^����vf{c���u��]��J�6"7�]�5�x��ĺ �5��!��{O�e����ʼsWNc����!�" �����	��Ɯ�SDPWu���w�EP�uT2#����s���$\L���n$Gm��֎CY�)������8^�z�>�BW3B���S�# H!�쵇�Uӂ�*�hB�Ā�j�U�9m谹�;b��4f��+�;����7J}�L����	���KE��y�x*�8��^"&���i���H_���R�v��pRh�X 7B�G1i1��������.��M�"�|����
�P�ň�7�6\�>w��B�(�X���z��7A5��VgO��ى^Z0ς�����e8-	�fX��>y@I~a�ݘ![�)��i
���*�=�����R����RBmi�kR��Cl�EP�$�p����8�J]A��EV�J�QC\�i.��jh�.?C��k��P����㢐/LnC�����Lg�� �� ]���4$IbX���g��˹<@)Ma�����$�e\�s�Y�M-LcU�h�A&������cɸ�"�@k�Jѿ"��C������~4���"�l95��"_Gi��J=M�����-�����>
}��wx��)��ꝓn���$ۨ�u
��G�ƶ���=&��w�U6:,Z��ŧ�R�G�����˲�i�cq�D�& �_<uf���r�g7����Q��4T+�P�L9���y{YZ4ὼwZR��6�M�oYڸ�H�����*?\�����j9�[S���E�B]���2V�)�!�2�wx��m�q5�o����\���j�Bw���ЙJ9摤^T��޺Mk��}/��$���RYh�A͙����r����#�r�:��@u�3<�K�mr��	��<�뛛x��*��8�d̐�u����ߕA�)�%j1��<�k��k_�=�y�|���q��^RRUm�]�[A�[���$��(��� �B��g�~�z�Lw?Q�.{]+`h�E{�n��H����ݓR�c3X�n��N;u�Ї�*��M��?O�acW'�e]���{��P!�{��e��]��Ô#֊�� �W�WS���v��2
����{�<U�����`���w���*��Z:	
`�fM+�s�y�\�0]eB��$���ky5S8�M"E�m[	��"���r�5�3��*�?{{q��o�|H���/���Y�YΏ��p� ��Uut0� �J���-���0h��L!�G�};H��m��)ۓw��yU�|�>Zy�A��-��f��I!����8�]������b2�`��
T�/��ϡ��Z@r��1���Wb���k�R�I�8S�(ns�������
����!L���k
��<�ÙZE_�Zxg�� ��[�(\
��cӰ�H��G�H����n:50}0�U���mRmT�*�oN�
��4�h/�����o�O���j6G���Yu7L�D�:�y@{�/O��Y�t-�+��X�=4��[�X٩z���ݐ����˟c���3��:�BN*�ئ���N��4c�1�\4��K�$�7u�gټ����b�5�K�)�n�l�&Ҕ��'��1?�$�1���0�̧�����0�WُP�����:-�鈸��Kiu���&�&���s���B�|\��h��i����
aRa"rj�+�,�h��x<o�PH�{_~����aҾ�����\��D�!�@ŰER�w/����?��y�t=.�zT�-���3��>��_��7�I߫��<#��U����`2��&��ȸD���v�*�L>�2\�QD�t�e�,�Ⲗ^2o�ZW��^���A5'��4���Go��;�����m�b=3�� �*s~��¹�����c;`ж�qʗ�F_M�+��}�z�G�6=�,��1�(�ee���A��_u�hV��U�t�%5J�T��5�|YĜ6�#�Z)W�󘘥x�� �!D�R���)g��j� 9�%W��7�~m ]-7�JWG�4t<��m&wD�ҹd�F�uP����&z6�����`�_�� ��	�l��w珖����(jv�]�Eԫd\j=�����]n`y�5�XB�%��F/�)�|2����������K��}<�ξm%�ul}��~�U��7�TLD�{ߢ3I�j׷X��5#'�ͮM�}v�S�M�
ٍcDd�4w���ˮ������Q��Ff�� ��i���( �H=+[�!��BS�Ͻ�D�MO�֏�U�tAl�!(�
�?�!�	G�#�R�
����%=�!ue}�nZ�=G���c�'ס�}��fѧ:�a�(��g�8���c������S��Vm�
�����:ߣ���9=��!��ͥ3�"8�|�\L+�(XԙL��ť�khD�v���^�1K ��9$f��5� �����;���d���׎Г3H.:	��.9�>�*��+Wg�$��#��GKդ���1�bTee}��N+?E�M��ܹ���e�(`:��D���8�d�`�����	l������Y'�ټ�MF&a>v��l5LU��I�v��m��<i�&��ǔ�߇�l�VǾ�R�Bi��Y^�;����,C"V�f,��Pig3����H(1�&���*���"K���U������G<Zg�U4+W�Gy�3z��|�2h�q���L��W��ׇɦ�a>"�����&d�,��w��aY��M�/�^tِ��\���YMÐ�ÉC�1)^�le}R��f�������4gU�Ԯ��_¡R����d|g�u&�Ŗ6����V�a��R.��&&bw���NS�>�|�곯 ;5�2�?.K�����+/��E�S4��b�ףc�����0�b(����^5��ۈ��$�fk�^��@�\e��@H���\���,���m�0�v³� �u�s/�s��������ݘ6T|���^GF}��ㆥt)^V6OCm��M;�A�?�h������|�B��@�u������P�w9��*oU��x���c<�ۏ�"[�JM�ļ|�LEٲ�DC��c�C�&|*	q�z��`4�����-��@r����}�R��ūaҭ�t.��v_Pㅺ�J��BY�-
��������R�3���Q����H 0i���8{zx��w"O<j�t����\�IN��RC�_�������ݴ7+�~�{M>Q�MMb]��]u����P@3x)���$�{5r���q����Xj��:7�Wm�����-&eN$p}��T�W��nT�?Q���`#�����/?�1��U�|��G�ؕ�>Y�V��Ņj^�ΐ�X'��%$�a��^���!Vr���ш(hi�cb� T���a���O�2 ��u�}�l:k#�pk*HI������� �Os���)F��S��4���&���پ��xL;�1�F���1�x�R.����4q��|��Q�d�i�3�$��벑���_7!���Tɠ
�z����TuQ�2?�92���\l��9�ֶu/��Ϸ}�B\eT���iM��Q*`4�*~6S?f�.��,�^E7���mP�*_e����Ga;�� D>GçĉO�[����n���jQȆ���<${�JJ���	��;�����G9��t��Zg�����$��^�d����V1 �b��xp�v�!�;�)���C�ph�v�λ�|Ԫ�&H�z ;eu��41q�Q�#+n�1��MeB-)���yx�}�+�$4s}��)�7��y��9��X�X���BJa���X�HZ#ԁ��J�O�)^��[F�XՈ+�e�R�ՂA�\�-B`q�e0& Τݢ=!U�F@�F�$�-�ڪU�ב���d����z�7����c��b����#�d�hަo��������{l�I���������� C5��F𡔄�����N�A^���y�g퐎$��Q�*�t!)�;U?��r�>����8P�z]��^�,^�p�B ���\ݐ�_8�O�׽7%��˙���F'/��(���[�$��
cO�]!��z�M�G�S~�K�`�����1��k���uQm���S�\33y�fS��b�vR�{���U�>�X�v������Z:$��3�Ijh�.����P�J�ʽ`�E!�Q�)�����]���?�&�}��n=*J�r#��Zp�K��L�{�H3���F%���qgj�܍����|�aK9���Mv�f���	~1g�zߴ��؎l
� �c4����N�#�W:�"��+#BX�}����J���o
������u6|��tKM�0�qbeC�	�J��ĥ8OP�n=,��lR7�U�"�vA�!l��Ye�7G'l:V�%�?d:)~X;�	��~){��B�Y����p��|�9T��r�^��Q�Y�N�ڣ�W_�(�F�]G/�9��؏(��̷ֳ��IsZ�F4`���)|`�Ԁd���&�e����Ƭ,
f�j9�Ύ�ˈ�2ۛ�q�q6���:�X���b�	BBB���@� �<�$S�5Ps���^\\<��+�t��N;$�9B�S贺�)��@Ic�5f�T��F<|�CȦ&�G�#��5z�7��υ��q�{����W��C Ω�f&��PS���Z�J!.�*u1<F�p����|/^^0�����bXt�|���O���"[���˾b�6(ɤsE�g���:y�����zIIK�����F�������WU]�mB�㖮k�!o]ݙ4��}s�fW�GL.�:�LN:fod�<\�Xv�t�q�ܟ�}	��X�����GJ��S�@��a{ԁ���^0����ĭN����:����Wf(ʳu��ه���};x�b�o������dM���V���R��~eQB�|v�"7w|o�_�o�`Uգ��2�*�n�̝����rQO�Pq�-���Sss�)�����,n����*�C �V�}��#٧~�c�C��+m�75��c��\�Um�����~�AW�3Uo��j��b�>�g3�x�D���;���^���NG��\x�P��5��b=IB��b�����#$�����h�E=#����r@�汋�����W���~"\���Y�7þ@$���W�r-2����%������O�E�_t��m��x��<f��͔��ֹ��dY�NQD�JN>�1��Y�B�����6�֟M�$�=jT��r�sd��AE��rz�zg�`�w��E|��rQ�B��➏||?L���O�C~	�krS_���z�}�2t���C�?��9hX�x�[����ozV�ZG�[<
m�t\���^�@Lm8_$[�.�8�x����������/�̰�8(F �*�:Qѕ����w�\0�j!�HGjTMP�5�9kU˕L��7��Y�UB�臉�d �k��<e����� e���̍�0e�J�:δ�IY����� nC�(�zC蹧�~s*���Z,�
̓R9�����VTDj۶uz�s�Z�C^����5bI�3
7�t]��T���w�	.$;���G7:�$��NTf~{h�8����������4E	�` ��H�c��^��t �Eft� ��4~w6(`+$&�\����k��K�EL@�������ۛ��ˍ1qq�g��B��i�u*�8 ���\��}�۷�9�~Ճ�H��::���N=�=/{���p��3>J7���d�r����hw(
��ZZ��G�@%�O�S.b�Y�i�֭}�$�-WCD+��ߤv1��ƻ�֣�m�|�T��v4���->�<c"���	�Θ��U4�Ta�S��`M��`�9��(䁘 ���(D,n!��> �)S�nR�gEZJ�|&��p��=Yb����nj���������sh�ȁЛ{�R������!9s�Eu�abbb�^�a?<��D���x$�N[
f��{��ykHYYY�s�����An�My���p~%L�0�\�'s	s��t5�z�x/u���0�}~` ���k<	:ۙ�1��\4��p��=�F���|�����y-���諸_=+4q�ЉG��; i�pMV�!��5��`�Le�|��~{ꦎ?s��|����z����`���(TbL$�
��s�c�|�X"��̀a����J!�e!���nT�NMM9�JI�v0�;l�*�_�N 23��'i^ׯ�~a�f�y�j|�N�
�y�䣬ʐ��^1�j(��;8 ���!���ݙ���p�~w�n;�y�םF''A�ӂO��Ff�� ;55<�u��֢1�.
���b�t�K���k���3���$�ͫBN-��S2�)����,25L6@�:X �\�9�Ez)$�N�݃�ccW("*Dm ��^j���TO��H��ч_�vPA�M��I��ڌ���A��z�P�9��^�3���xT��;����=BAA��������\$�>d������d�fi֛5�ԙ�R�7,� 6]dյ���^�;6+j�B���R�|�2j[�T?�1ax+��(�\+��~�8�5���ժ�ުYr�$y�?t *!%�+9_	CUˏ��I
::�
�{��q����,b��4ޞ�~;s�Q����)�Q�������|ZŴ�-q�z��W���W�Hl����t��2 �<�o���`/Y������ ���/��b���4-���))	���4�X�)/��S7�_)R���Cb�F�9b��4#�u�B&1����IG��'�S:��	: �0�k���*�m��e���ᾟ
q������׷)r����ƛ����p*��qG�4,5��U����(����?��' tc�����6.�I��Y����B�m�5�M�(*b�98�/U��?������`��Hi?o��/��=0/����Q��St���j�Ge�m�R����P��򧚱�Ώg֗W�`2S�\�z�
����������|���@~��G��'��~��R��wH3B+��;��ʾZ*����~9�c����s�P����g���.'DZ5�t�d�naa��H��h*�W&�-��B|���|�����Ŗ�)��C��˅�4t]Z��Ў�-M��k��۽����Ǩ$9H"��cQJ��~�;����x���zk�&u��U�}:�zû���}c����������b�4H�_^ ��Ǝ��og��/,0�)�H��{�����I_tӎ/����NJREh�c	l�|rŰ��"�B?��K��v�.�@�ot�D�h�eee��T}TU]�6
��HwwJJ7"�Hw�t�t�t�tJKwwwK׿�������z���Z뉹��h�v܎� �wH��{O0?�L�!J����z�!�HR�gl�T�&jZ�_�#���@y2�l����o�tc\@�ظʉ6���=���17>�K����,�|���1R4~�;���:6#C�UX�*jj<ey,���<
�W��J9�5o�b�'��0L@�%,g��Ȋ��	`�����w�Q��;x(k��s�O����u�J��P"=XW�>��_��T��u��L �|JWsլ�:�:�b�����D�����̖<�n)���,R��ۭ��C���4@.&����ϯ�'gs�[����m��&n���z�dh9f�`@!g�ghW�k��^�a
�T�>��i4���+��HZ?X<�h�ѻs�X�� � �&m?)R�ٸ+��R��'�����! �&}��z�5��ji3u`���a2J�������P��KDЄC���(l���r�}x�p��\ ���goA ^;��!	̩����!�� �D�A���SW*jj��Z����W�����zt��!a�ӿ����}�f[�����nHK�q��]:^iD*]-��Q��"����t�<����\B���WGr��T��)�k�ZO�~X���,��u�L�^h�y�b��Y��M��A"�uTՍ\��<!AD0a,�a�����:0wG���߈W�ښa/Ӄ��������T���#O��Y��D�N�+����y͸;¹���fE����1h��=���������"k��s������&���f � ��?B��˾����h��q���/ǌ��[D�s#����i���4AN�����^�K2��p[46V������->(� �?7��,�����X�}<��G�r���Oܞ;#��1h�J���W@�F-�t-��@lvs̆g��Ԯ|�)�{@��O�L�v0�:Jw�����Ą�I'��Q�F	��ں��,������?�ׅ�3��[-�'���f`m�ѽM+U*Y����ݤ$e/�DmXXx�
,����!y��S�����M�C�ɣ*(���!h�����w�ih}��� *��b�3`����yы�TA ��.�(�l!�$4��O�v��ղ�|A�?`JZ�6������$tئ�&�c�өK�O��v���rS����E!����������F�gNz����Lϐ [��e��'�,Xf�s�%��4�����Q�%Ψ��dfʥ��e@��R,jQ]���!i��!}����&K`"!x�)��xhhh`` ����olW_p�V��]�(�l|kAJ��J����=�r�����/��-ߦ�~Yĝ$�mEr^*���9Z��ȷ��w������]�'\��z�|�\�q'���`��@q�� @:�v[_�Z�Fy�~�� 0��x���CN��o�h��0��/_�Ė������!0��(�l��/n�^�ކI�����5dl�m�~�TQyH��n� �q����Tt�fXKII)��� 1%e ���/�aC�T�p�`��`���N�o9r��2�'�ù|��u��|����7~B�M=��;�:f�������{�#8,:=�Ƞ&��|�mP�U�9����|#�����K��xtU��g�G&�f�ߎ��8��֙�]��&+�[��-�MFRU53�;'/�2��)�48(b:�բ(�qFGw��� ���}��R��bm(0��|���i?��R	���B��<�o08<����6�������x6L5FъJ8ݮ� f5;����ܠ?�Xe�(�<c;�a8�ww>�i�~wG[�څĹ<~�1a�`��j̴;I�����S_4���7�� ��V�v8�qX��H���v�R����ܫ�?��g�s��A���м(5��r���o�Ǜ���w`��"k�4��uݖ˶eE�� �����/1@�y����G�zn �r��	v��|�lGgU�\?�8R�#��Y����鴥�Y�]nEn^ݧ�f��8��f�w1[/s��y�]�2{�L)��6t�ϹO�����AC��0�(����\�jH��X5�h�8r��f(}�x��`�Ւ���ƀ����r�j�L��*�u۵���m���o�(�
���xj	����EmٲEΛ,/hg�pj��?1�K��׳�b���C^�ӥ��`��
<��\0P��=8�/��ol�<]lh�\�[Lq9���y����"�{�z�Iږ#O
�&̀C3Ԙk� ��=v�#�wp8Xiq��G�)Kg��ӤS�����X�������;�G#�0}��J"T�����1j|}y��<=�y��s�M�s{8(�	w��(�͑���������l��@.M�[�?k�^Ֆ��N!t.��%o�{��O�/�6���_�ò���2����3���5m,������F�_���1Ŗ�b,u�pS�}��������I�����ũ�o��tɝ=I[F��cJ49�M³n����}�G­Xi�P��ٴ�^Tv��
�^���b���q�������c�g��lS�����{`Zc�}R�f��]�=X!m�vբG�˒*Γ�/�87Q�����tGz��-ب5����K�3�WQ�@��������AN������
/@+QG��F37~���!u���ƥ�V�v��z�bh=�r������������?�/����_�����i�ܽ	>��m�W�ۇ�����^�����qɤ]<d7�N�N�{EC�����I�?< �9	p_�Аʯm�H�䀍�1����mJA��+@7�zJ<�0W�� l�]���24	/���-����Ik�O���D���C��͉���`�vd���ƈ��M@B[]s�El����w��ڶZԏ����c 2�n��L���������J���z$��M�~��f@����R0��ە�3 %��~x
�HC#5�.A�Җq}1�`���@KK[\Vqt'�'5���$m�3���[���&F��=�����S?��'�VJG��(��(��p��Z<c돒B�;}��.6Yhd|�)p��v�;�n�������e�1�"��M��&J��|AcA=�C$����T9�lY�����n|RR!S�,��^k�^�:g�-xV��Q�~�c�㧡�B�5���E� w�aJ��b�>��Rbq!�g��;�56_mx p�̖��b���>�h��BґY�ʐ	��T�T`�ɁRi5`c�U�|�k�HJJ���f�>�� ��*�I��y��ḿ�cR�g�{H���T�[��Q����yv�#B����M�O��k۔΀�ޜ��x$n/`64���&ep.�~��)T����H2����6���\�-o�	Ъ��ME�S?%�M0N����l\N�?䫴�6�o6�|�?x�זO(�����l�-�� �I��k
Hy�uPo���)��r�JE��Id�s�?WI8'�ˇ�Cs�� ���}�?A�>*�շ��=���0�
���\���60�9mt&w1���?�8%~H<��sdخ�2S�h����i���}��Rd�3� �jP4��&�����҈N�9�0� ە��[hk�o���P,C�
�j9fl\��q�Ô�R��U���2�����\b�zޡ�~ zJ,��w��]�&��4�?7�7���e,s��T��~i���h��0�c]�v�LF]f��G��[^}�sp�AV������̅8�h/��p��*�o00X#�@��_b-�''�u�X��irأ��&�@��o����;c�fŁ�0Xr>�I�>>�<��$�����W��P��1O�CF�_�V�4�mi��Z�N'�Ve?~{KA���yP1�[��,R�3�V��Ȏ,F��!4��s�bk:�2_�m��V�;�Na��w�Q.���2�)��'����=�dr����u��C�]R-F��6A��74�Y��KK%Wn߇����@��������`����=�}��|WZ�L ���0G�e������-�^w�Ϭ\ٻlw�4k�����0�=��bV�lc�z��l���.����,� v��/�
�:�=�=���'"��}Ԃ����:�A�C��z>���W$C�g���9"���!�5m��;���y<X�D���+��F�nW��s΀���Md�ц�Q���BF4�aJ�J*j���.���c|W��.�P�/�*�,�� 7��V�p=�@��J�𦥤�7��LO���V�)���S��A0���!S��V��延��+(~����8�I���	"�JLH ;C@pX/'��'@���Z Ӡ��zMq��j�������ѿ/��|�o����k�mK@(����x���Qma�t�Y�� �զ�8��t��� E���HN���I�ʻ��M쎻w���*'�3 4�ğ����"S�۾#�?�8�����u�O~Q�E`zY(ނ!a4	|�3���^�hM`�]R�+���i8���N��=�<�Q��噎eJFv�¬�����%��O��M%��ջgB�MY{ �r�m�U�k�Qr4�5.e��G�v�i��ÍJxJݐ�и��`Mk3�����pJ*��lt�v���w��p�-�U�#��rM	33j����ˮ��@���ZC��f�B;��1gPA(
i�g�u��LFv�S@tπ{=:�����x�K�6铓J���&���<$`覀�������'C�f(�ҵ�&��L��B�yB�����8܀���:/Y�����{�("R�-@g|�1���I2���kS{H͠��.��rH��ɱ䢧�O������tp��<3��a�U���s�2Ə�~5|rACfV��	��5�fW�u��%0יT�v�4~<*՟HyS����a�R��E��Z�w����ԼL���,od%���
��p{��D��'�(Z35�ww�#�t��Op��Ŭ=�����=��������;������d��K4���`���g񔵴�(��	�D@��V4��* ��P��ĭ?m&�$eRي���I^�:쁥T��xc@'<��������[���ۥX���cl/����\�eK����ʬ�����70�k��C8�.����U��%����<yHL:M6�����ޟ;*�(�x$ `���EهPV�ϴ�������?��~��~عx䍦\�_ �Orx����٣��(�t���CX�/�^�P� �[��(��u���5�!�@�4�[��_�����a��42��o�&(Û٪�2�ݯ���a�M:.5�t�=.�E�Gf���X����Iln$�B��77�ƬzSNH�K��b��G�`���`2�+p�-u�-���5X?Ǵ�hb�K.(O���|ntZ��A�|�h ���B�����d~����4��X�_�c&��nZ^�3`Sr`��,5X�
�\� ��eyT������x�3�uᲅ�o,ZT����s/NVʧ�9�Srҋ�333���N㬜�Y����� ���f�\7�+D���X������,;�e�Q��4���q���qrgUڏ1�`�6w��NY3��p#����Ay����g������wʶ�o��e�Mx���8CNe�6��Q,{��ɹ�dkb�d"���^:{�:Q���,vӖ�K;Y�g����FM5\��%���Ү�xI0��y5��4��&t��c��L�Z�^���Vm���#�U�C�
���3CH �����t|7����Gs�p�w��|d���@���/v�tk �Y��.,z�O%�Q�5 ÒYM�4��p��{";5-���@��]qѹݎ����j����#�AGM�Xx��E&�q�!*�	��XD�Pa��]=��G@�tz��E���p9v���E�@�纉�q>F:yAC;�!�Q� a�:Q��N�9�廞V~:��!�4w�Ԑ����h���k����H��v{���X�%��¬�-�̬�GBc���7��g"���и�y`2�p^�E�]��6G�V�۵jCP}�<.����)��M��ݶc$�����\|��p�-Jt��ج���+�b쮷Dd�c���+A��֯ �l<<�Xax��-�U���V�Bk��!��d8[����ET�8J5"��j��5,}
�m�z��aOHx��/�>��s����5���}~^�3�=$���}�v]�"m%�����|�� �R�ug�'��S޲�H�;θ�6�44L���ͻU��"'��ٯ��Vu3���%3u���a�:\��a�,��Fgm³g(4�p������WƼl`����Z�{��>�(��W- 2��y��a�$�XA���q*�^�� �P�r���J��@�Zd}��O!)�˔֏�b�qn�G�&�w���!QQAB�
�;�Q±軲|^�tuu�R�o�9�L����Pd�S��^;?�B�j�g� �X0�R`�F�:3!��c�$�䐙i��������Z��X��<J��_`4�p릛�hG�ͷ"�S#��$�8��Wț�U5:{SJ���7'�Ą�����d�<�<��;%/uS��"?!��=���כ׹ԍh�|fA}�F��
]�5&j�T�h�}9	�1efC��kQ�?܉&U��+#حѝ!t ��C��S����t�),$�cY)"_&�~ä��'B%�Wڽ]�R�W�Y�"���-}Ƭ�v�!TQ	q�� �2�ȉ��p�FgVdvv+M_MM�nZ���|��r:�_�~�nZM49�6E���v��q�]l�-��)�K�p�q�{� Z�&,�w >�{���R]��c�F����VKZ`6�
���0T;j�אڲA�G{�c��ឰl��]�� �������g�����1��G�����uY�HTq�)*Ǉ���:���<ل{0ob���IS���F"�c@C��f/ ��)��p�.$l@BEF ���I%�;�k���c��ǔ�����H_�#w2s;�*��^�Mvn3a�-�x��$�#����9n��hW͂���q�]Y��/`��d�a
L�|�oA��d9������" ��A��!������V����ZƙԞ�.؟�s����>�ӻ-Q�'s1q_&-��**���!���`�O�sp԰ƈ]3��HE�{g(	kvמ����̯��� � M+��`ѓy����y���b�Wn]̻Q��E%�^,���-)�4�N���)���6��o��=J�����NIPo9h��A-�;�W��D)O�����{�4E��Pfzq��}y����7�&'�N
����o�M	\�Ș!��F�h���O�n�VV 6S(��e//w�4����c�&�wR�%떯�?;�A���?;�r�����Mh�<��d�j��f�|���b���ă���gf�����������M;-l@�QQS�555?23�jk���ȈIH�89��ܑ��R�щ��d6w�7;͞b�{�557daQZ�G��W�؞��`��������/���&ɵ�ᢉվ�>�
�L�ё��z��^/nr���(26��^�ǣ�ĕe6{ѿ��2�]{CY��'z�ң�������ҾOвD��wz��f�-_7��Ê;��3V�?�N&�Wm��$�D-�eν�2���v�l�����&� �	��g'�Q���p�t�T�4;�De���.������g�~ee����2~�����Θ��W~��~�/�j���<�������;�a~~��a�H��NL�*+/׷���	����F	DEE�����d���������×bP�&�a<�} \��G8���>6�#5�.��2��}1U	s���g1Il���ث֑�5�^�p`C��2As"~yyQ"�j�����l�����ȋ���3G�N[XUSOO����p0<��9�a_Dg_$*j����T�Gw\.���w�$Q��t��b���)�ѥw�
k��iX�+�z��OE�h%>9���'K3���SX��FM:���*��x��<ɞn�Cg�c����f��1�(��E���|`ҝ��?�$w
iL��b�s�LoK�����`������NAZ��B�g�=z�*�t�|cKS��t�",,���������ol��ﴛ;���@���F�O)�qU�A���k�1.]|�ؓ�+(�a��u����A`2�u��В�m�M6pP1Vvb��=��p��h�r� I����8���69Uo�lj��6x���N��� p�ϒ��.�#4 #��C`�����,q�D�Ǔ��%�|L�K�8'��x�˖��6�t���솛dc3>ٖ�)ݸ��G��J����L�,/�Н�b�=HU������x�cj�c�"�j'|�y�Ʌ�����\�K6�o��G%�7��=����,Lll=�q��2w��ui�--��++ն��33O�W\���:�w�Q���'��F�6��hyQ��zJy1��])(^�>�T������?���������r����C���K�������_3�`��/�.�˝7'K�����p����i�眙�P�R�AP�z'�������,�z���n��[!)��Pjp[3Kj����A���n�IJ=���,6�5��nH�n$m\�ڙ��>���0ӇTV����v��CIO>�VלDi�lt���YZJ���j�~0^��n��&�A��6җ'�d6Ifdb�9�#�e����Y|:�"�eMe�䏬���
	*n�@^�PG�x�&�}�3ְ�@v��~��k]��|��Xl���ɍ��_Uu�'{dtT��������!��kOB◜��M�x޴�3i�w�E�{�#��#�ha�b��(`?�Ob�;�3����k��2�aő\�_����p<I�(��,=y�uT!j1T^���"����/M~cKNK��\�莊��EA��i=j�GǠ����������H���rS3�>e<Ӄn����&���+�jQ^�U�\DP\��K#��ͧ���r�K�H���KVi�J�2ǲ�Žn����v�������+�H3%z@��]@��`C��/]�f{�����ۻ���64�Δ�nj��b��pܡ��J�	��_x1v8x���ZZ�$F]��Ya��ts���=Z�]�	�E%�40���Q���#ml8�6���SU�\�(�p�F
CH��������m�DGG��|<�P�+"�R"�7.J�Wwy��=@�u{l���s�=W�(*+O�������n�U�Ka��^F]�0~bS�*���q{ۊ��ǼQK2_�G�'�XA@�[�iT2����F-�DO;��v�-�;T��~�D�5k1�eN�i#��4i���{��浿q��{"�s��"BC***�O���u��5E��m�r�wx�
x��<����"�Nk�}�:��T��,r���L�$PS05�T��n2��1�Ȝ_�=]d��s`�#EV�nR�o������隝R"��N{�6����B/�ܷ�~:܄�^H(x�f$�
7h�A���o?�^N�b.
����|�4K2�fU$ppp!��RR�SS1� ����{%K𘘝
�����34����������B���YՐ�D� �b�Q�m�>�C��Q��4'$�/++��z�GYϬ@�tK�o�1��eeO�<D�<����d�u�[|�b�w�q����ҿ���f��_Q���(����ʂ�������J�z��m��)oS���tw(%&>	Rtwe�KXe��TŖ����Q�v0��R``�����|�߶�m�u�,ŝɎJ]��R�k��]�����p�Sع��"�ﲡO�.�'-�K����8�2�ke\\_���7���pS�\�;���6�l���# �O�
~����Rwl2�o䵐�����L�¯]F�i=�h�&<��݁�/�F���O>ƋI�R+	@@�8�`��R�r�����%��v�7'}��[�����^��������
[ZZ�=SPP�p��}�TG�-����̆L&�8Z��je?\���ٰ3>�&L>2�7�Ѱ�V�F?<�{>��Ί��q����$$I��g�?�b�e�N�>H���b���&�R��,XUt���~N��o�D	�)��MNN��z����#/읞a��EM-
��F7R�K�T�M�l��syw��q~��>���8��EE)�����'l�� �-V�������p�6VT:���=3=r1~lrv�j
�-�����u�����*��k����h\�j��)R��̗�~4_�2S � 4�T��Y'ԧ??�O=7��@	�n�)�����ǳ�����v��j)������OlD'�?�2�Lo����.�&	x0Q�zF3x/F8ײs�o�P�>�
�%�q+�=��sE�~�M�P* ���"���������?W�}���ol��eק;f���c���f����R&���8�U[W�P��J|A�"�@�9��Чn\��P�������%?�|���;��-��&V�����|D��.4����B�

�.���L+�sw�p����� ܄�f�~����s�#-�[����C#ø��N��of��0�oN�^��~_Ϝ�U��\�V�;fzq��6�bF�����x
"�zW�F��U���	�̰��6>�5wjT���*0�[��	��'����!XH�jo������>������h.����ݻw�pp�>�EDDd�^�Nf�	F��H�Ɔ�Ƞ6Gi�3� (����İ~�!7�,,����-����Z���PV;�H��!5X��hg�ݏi��r��L{2�W����7lã|�w��'GMu�彿;��V�?�kL~6�oI^6�Զ�V�چĒ&mGgg6�ce�)E}��f�i�@��1�Yn�hp`�X�`O�>�ƞ�7�"5%�x�X�:p��b�C(�H�H2jo���e���fy���gV-ԫм���������@�憁�K�nV�ӏ�<��'B������i8��	�R�i85U�?3q9c_�}	�T~2�2���G��+�{�
���\8��g0U [Nh�������j��끭qy63W�T�_=��k5�o|�P$��==t�tm-�޸ �r��Q�	����Eu>}��RTPGFnh_�RUQY_���r='�q9��|�8�.\�����n���A��ި������Y��Oo
䳢�v��i`⬏S���Ҷ�`N����3�lV�BNei�
Bű�O�:G�����08��ۅ�"��v*2����Fvt�4V�T�ՠ�E�ܓ�7����ON6�cy�#5���� ���8�=%�k$� e6�����nk:���+ˊ�*��#K��5��E�J34�k��R����)��:���z��0� f3&��M�#�������i���w���s�ooi�֒�-�����T�3��|)-�m��YcK\[�.�#5����%^ws�1x"ʊ���Â��v.7F 1�}�R@Kf&����LG����r�? 5�����z1aڷ=�e����4@д��*|̭mť6ss�`���QT'�*q���m��D�|}���ۊ,������@6�Y�������Ն��i߈���HQg[G�>��� �"�K��qUm����h����Q^��d���]���.�7o��ǁ�~�7,�|e���;{J�4?|U��Р��g��D>�T_�A���	s⎪־9����79�$Gx�������Ĳ[r������\��.BE�8��<VA�qqteC�Y�El8Fi�3;�����x=���ό�I�׶7�B���Hy�P�0?VVa	���PX�����L$�P<�3$\�=S$4�WT�{�!����ٜ�]����g��	�ɺ�����$���W�{uK��G���}�i��?��O[�`�_B�����F���:ٶ���w�٪�ɲ^8?���ۛ�>� �onN,���z>�44�]��:ADr���I�lk_�Q�*����t��ʏ��H[)�N�!��k/{�����/|��%��������3�߽���.�d�*�'A���!��iL����x(��)#�w�<P�ﱰ���Eȓ5Ry�S:�Jy�E�G~����0���Pe �%�e��$��\�n[��C��a��)8�QEJ���}5�Y�`^��n�����^�v�>(.��8Zm�(kn1Ԟ%��S�U6�4/79�y����%G$XJ����Ε��n��k�h��z�x]������T�Y����	{
2����RI	؁���a�݋7@����
>�^3���k`@��Mb\���\����Ͽ;�rBx
 V*S���17��ۀaC����?�j�Y�2�n 8����*ժ�
�F�2����X�f��ΐ�8㕴�'%Q/ބ�WB&�h��Բ���5�\��8`g���O���a&&&\oW\�>|(>�&VY&��$��&&&1[m����^�M�=8<�T`���}E�/�D�߰|��{�<��5x*�8�3�<[��߳|��f�
F�����a����g��l
�|�5�FEG����c_b���v��Ѹ��QGMYvN����HM�������R�y�]�������r$��� ����Y/�GFLZ�V��r���¯�,���"*Q1����do�֚����iU\���a]Y�000���q�F%juC%�V�1'4��~��� h� %ж�3��#��]`����!:!mm�y�w#��[7%���ʇ/=&Q��1H�����p�[]S���E���ӭ�N+��>Y�O_���	��_�5�尋����f�?N��wB���ܪF^>:2��!G7�![iI;!+%e��vS�8Py����b켷@V�H')�D4a�_�z��-9�2�BAr��=U��U�I��L���cH;\��妓���8�̖��Iu��9���;W���V?�����G��O-"��u�<֢�tC.KJx�Z���E��I�+�ޢ5d~�������j�������E�����Hqb,���Ş���B�Ԃ�^�u����Wx��c{8����
�t���+�e�"���G=K2�p.������KK��i�v�z����,o@ >���a2S3Qmy��,E�C2���s�`����Ȁq�pllm��{�31)��"�2(2	�p�~Ep~?$���'�BE��i5^��ۏOj�Z�j�sý��iq�~�S�	7�?�(�X�(1��F��F�j�6U��H���+�l��lmm��`͞f�)����b��x�b�0�3�����K3@��Ĕ��B�)�c���Iay'�H�&��m��\�u�(���G����t�8�S�H�zMҸ���W��"���D�S@�4�^|���ʫ	�}w��F!���E��G�g�[����}6\q��O(��p���U���B�2x����z�4A���0�*�'T)w\ߚM:��y��5	�~���]@M���v���|#k���7�����R:�<�!��і*
�������Wt���w���	��=g�����L����{xXf���b D�����fP^\ѻ����\ЏS(_��X���' �T���/����*��'�H�j�F����H�0��hzf̽7b�kkD)))���J�\�wLA(Da
p~���4����C��|n5��x��=�b�Ę���7�ݔD�^����v��;g��BON�/O��gѵl�d�2�666r����U]`����B
|		�)lf� }P8�v�À13����8��b)f�x��������t��x����w�!���q[����ܖ�{8����Z���U̍qb��
s���=T�GR�)������Mp�Vʂ���놅���NK+9������]X�Z4������g�mJ�Y�X�2�Lf�,������#�Q�Q4��<7�1Q��Fp4�� ��;^�Q8mVrr�㶴���=n�Q)���QZR+O���W���"�!r��9�tW���0y�������FL�`�`�"���|��� ���:6���������dB.(���z()Yz	%��J�C#%��b~8a!�ҁU�F��b�h�F��
t�o}����'���L!��X���iT�I뮯k��,W���>��\���b��@铴t逝r�\��P�@zp���D�A$,>}�ۀ�$9����3�3�|���`���]���#�w�����T+FL8���EG��^w<������}����j#B^ъ<��3����������4-�����
*�:�<�p9��ҽ����:6�c}��15�V��d�=:�U���ƑK�?2��x��*l����/�ߣ`�܈���6}��ES��&��������
��˵nB�h���^�?��0N�Gvm����n�r�ZT,�v���پq�-3Qu{7)#����ى�h���|-F>b���'��n����se:���aU�R�Ɨ����>��z*�r�k@����E�]�s�KH�HD��FGG����+�-%��k���f�F�Q�����`������E*T�}�XJG\�{�C�&SiPr����v"cV�n��ͩ�����B��$����l���K�ӳ�x�_k��ܯ�\��]΢������3X)�ѯ�����,�h�X)Bf��n�M��7NO�VZ\��0ppBȥ��sD`�������R����\7tJ���� cnnm]UvԷ|��"�셼.�ϼ2,��7�ж�FP�b+1�:b�0cJR�j:0�V�z9��U��8�)*����#�A���C���.��H���3���0^��H/��"�Sp��p옲�M$��P�N�o�r��,�UuO�`&����w�I�T �g+�F7'�}�W����0��?,.AES.�dN=H��4n�9�	�[�x�Nˮ���\Z����������p^h,�ԛ$�[QQI��M�O�SR�⿭$�bC�z�6��^��;7;;[���%�|i�A��^'Ve�L.�������;�\��bB~w(~�6�~P1����������/�I��D�Z��A�_?���t��T��{������U+�<�*��ॉRox�'CK�ptZ/�[����_Y�����l��w<_I���R�F^60��_~�1��Wn��������+(��a�Z�#~����j�F���,���@!���C�������)�	j5-��'��x�������3mk8U�Ü��y���I);4,y3�zQ��9{L�R�����ܸ�HL1t�_��Fr�m���M����Lo�6�f""y:��&A�Z��݈V����Q���=<��5d-���b����N��5_>f�k觧������جP�'��pQİu�R]+33�|^�z����eӿ�13���y�kk��ze���ܝ��_�N�9^膬��6�]+̷|������Υ'*$����h�4��X�x��t=�+�xtp�4[�q��?{����Q�Ȉ��]���^�޾��F����Z�%���V�Օ�B.=�E,���n��ǿ�|����lǆ�����Th��]\\��)��%tJ [��P)����h���<_�D��*�7ʋtτ���	���8�ґa�����+n"�FJd�՟�ҹ7>3�1�]8�6xHBM�y3�DG-����p֤�l)�'���>�����`���Nf�!1ssB�m��Tiu�5�n�"^�&��������٥�~Y�e�H�F��j��I�W�'r���;υ��M��%��e��:��=�(�0<]�ZD*����g\��H�27F�-�j�ʆ�]���tޫYE��[Fn��@b`h��	cb���Q8�{x0s�9/Ez�F�S�^�i�3��?�������~ �$L��3ɌV*�)~�>���n�=ug�����ײ�Y�][�RT^*�.Μ)0�WcS��u��|A��,� OM��n����L�"�X*jjaVi���t���P�~���e��h���o����*�`�߭��N��L�a�T�����-��r�b�S��k[��:;;��@͹��>36���juUT$�:`�1]���y���0*��AҼ� bw8�?����L��z�#5��������8�'sXiִ��!���㕡�������1���ur�=����m�Rէ�q�䀷��ݥ�}���&&�RaE�[mn�F��['|�լq����^'��U�Fo�71)����t��-�)��/�i`@�5�E�aS"��8u6�G�m��ՠr���Z�9��U���[ZE0y�0�*�O���{���<�>F ��Ϭ(�NԏD�G����-[�w�g�1�<Z�Z��:��Cח�}>S ����[Ugɓ�Ԇ+v���䚪��m}~�EǱ��F���K�"�U��_������%��o��%��f�&r_ԡo��eύ�3�H��\��-w.a��s�~/qd�o\��(vMk�N=��i��Z�,��c#_o�[:���#�����1����F��Q�LJ�C�n�|}�"08�i�E(���wJ0��u)�\CKm��oC���5�[i��R��;G���Ӎܪ�/j3���I�^�}r�N%d0�M��T���̾�DVX׷�����}�JZ�=�8=�����b�7$<2n��~�����1bT�	pq��w�RB�=?\��8[�J9`bamN���yܢ����X�n!�騊��n=�*�)
!wwh��؏1�،: ���v�G��X��jC%%�x��.�-a}���tt_��X���A�+r.y��9�B�˞���s�u5a=�}�	�E=O�IW�:"���^��3$W�����ߏ��n�t{!���j/F���
�ͺ�|�n':F�hI��7�����o��֯�%��f{�����:ս׮�9%FϠ,�������ҝ�<&�+�ږ	#YA���Y#���_^��
��U�8���k$.U�g^����搪�6�C��^�ί2Q�O�`|���\/�2W�i��V�a,鼫�u���Q��a�M�َzKTH�t�`�_���&����m`uLT�%F�uW��"�3	���G�[�U�D�Û������.���i)I	)AZ��A:�S:�A�w�s�����|`�'f�o̬Y���5�w���5V����O54����<�%�ݓ(��bR�v{�<����g,����QKvvv?
y�����b�s�ܬ,�S
�	����c��,,�������q;�R��{�����<�7	���ܺ]�R�X`�3���a��ɕ�Q�`ɻ9��������ZK8��(�ꀿ��52Y��h"h�\��������P>��~vvD�m9 ��QS��^��u�;���k�B��&ИZ���Loޡ8��c�	����a�����C4y���񗳋����jq��
͐�2)ё�V�/K�������C?����-�k��a�g�~����*�y��A����h�gy�v�G��9��,?�����W��4��)l�S����!��Ah�o��L�J��&��FQ(qjx�0��t�����cmn��G�/���-�1C������o_��T�R}r,�������x����/Z|��&��!=m	jr��RC�D��i�{�_R{aR���9�hĔ�O�juu]s��%UV�`bRN2�ImN�j(�}M�FK3!+�B���&�_-J�H�P�J��R���[(iN�¡���_�����}�h�mVs$�UC��vQM �

I��F3xs�o<��9)��:�9bWǿؼ� � ��ml�TrDѣ�(o����d�((*ڜ.Q�#����I\�D��n&��l���T��F����G����^X���K\�.��J� \�|��vf*9BUghs	�q����~������&�jx 8�uF[��TC��ߺ��h�ŝ����������6<X)���Wx���ߏ�LʦK�^��r^!*�gA�h@�,i�[qZ;{�J�[
~��L�e����{	8a=�o;��UU��!����4�>���lh�pO1�r��M��0�jǈ*!��s7�m$������a�!���x�4>�.�d�6���Cv���<ݜ�UgN��H�_"/sf����$�`�+��f�I�X���̬������M�:>>&�w|���J��;;;Ɯd��"�o������
����pJm����̴���wt��\C)�D)�Mޯ�xG0��'��M<K�yS�5ݚJ>���#�[�Pg���=C�7�w�N�&=Bo,oF���K��s�����1��T�ZC��Uo�v�bﴬo�	NO�fޖ`!�SrEG�O1b�Y��n��m���ؾ�"�}�^��mdTyn�P1���H�Ȉ��/�J��͙ށ�k�YʯÇ��pR�
��ۖ-���j�-�z_��ԗ�d�?������k{�n%�L.�+��zY�s
��\��mM��ۈn�Q��E�=[���g����@7�2���(���2��ٿ�b�W�W���G��ЄCƃ��,���eS���(D\f��]�$z�s����/��>��Χ����k�"��?'L�K�rcS���ڜy�
]�<�?��E�B�@�N��	������wu~� WR\��BXW��1�3��W���uqz�lS󟞆��Ɵ0��,������Ǹ�t����T�'�k+������qjV�z�x73�KaFF�Y��,��qb�ק���ιzs�%~#��J� ���,�L�����3�YcF�Q��o+��9�gL�r6_I������%����w��Ԍ��;V��^$�|U{�;U�D�>��^r$����F��fƎc�ދ�v��f������w�8۹�ȸq�+��K���z�}����e|�<����-ډ�]��V*p����U��x��{I����X�`�퀊�b �ҕ�Q���8����7ӓ_�ي
�b������U�~��8ZXX�>͝o0	i3���an�,(��S�q?a�����V�c�G9_I2�/�0�;>9�*!z���}HHf��D>
dЁxj�NF�MH7�iC�x�M1R-<w�eMI��Ku2]�4}n���ֽ�p�	%hrRf}1�G�򵅅E��P�L���8%&&����
���\{�j��PA==vp�$��[}���*$k�G*�f7Z����Ʉm!8��W^���0�
[�0�~��樐?��-��o�*M��T8��Y�-:3������A�6FHx}�2&F��7�qz�]$�x��P�3?���B�� �/L��t����n%x�o~iy���|��1+fH�|�2B�r�Q��5&�X���9|iN����I�8��V�3���	
�SC�Qb�7]\���>�{��Q˞_�(���Q��%(C+���֏�7Y�PXn���tn~����(�u�x!�v!_���{x�����W(�ty��W�������S��� �D��� MR�y��~�\W0�	C�;�&��K�D���E5�[��=������M.��o��OV([Z�襓�x]�H`�SE*p<��j%��w��F=�wz�C��g�)Y�?_������OYk�4'Yx�0���5���K�p��v�L&�0��F�:w�m�aRcR���p�A�i �c��;JI.���^����%۹�x�"6�<��TLb��ޅ�&��j5S� �I����%�~$鍇t5+�P��}�D2�	����&n6�:�F悑W����o�Q ��ǈBє���e�QO�������5����LX����~�ެ�c&zO��B{�d5���L�RN��h��atu���F��W�2��7=��FN ��?U�k��9�&f�t�|�����øZ'O����P(���������޿�*P;�xXPFYo_�����a�`P�0)~,Ñ����!�9�=6�!�+�����y��7�Q�P}���ccF���Şg�7I��Ԫ��{|�3�9��tM��T�y{&�˿KD�|H��LIQ�I̍��З�~�:A���b-58$��_ [�e��ò�Ĭ�Ak��T^^�x��u��tSgzzz��b����.[x�r�w���FW:喡u����K�����t�0)��$�pa��膅[���KEﮍ�8��"z�׀�_K��VD������ns��G41�� 	��Ϩd���J�ςn�@����B]��)+&��գS�����_�m�_�~�	u�������?�Y��,R���	��7�pqr2Q覩�*���lq:
Yȗ����s��
qsD��~�D�wz*ay�eO���:U�r�FFFM�ͼ���1%�qs��_WG���k׹zF�(�9��0�=g/���tn��Z��w\~%!�!��)&=#�{l[2�k ����x��;��L:�X��ɓ���Of�q�U55�%�EP%��+m~P���?��E�L�LPQQa���;�����*�jK��c��.&;[q��Ƿ
���l�P�S\�$#K_(T�!x]���.x�Z������h�)չ���s ��Tӄ<Xg��3��0���U:y�8�' $���#jt����6����P)3|"_&�n���6T��������'44������ǻ����� OOO�h1A�E^A���Ԙ�'f2|�h_����bQ���`��B���"/�T)Ԧ"��˩��/�����ǧ��|������5g����]��bf���D;'�}M[{{�\s�6�2�����R�9�ƒ'XV��+(I�Z:z$�ϝ�����2B!L��dC{"p̎���E߮�y���$�+W
x�������7p��8�=����(�-�� ���Z��rݐ�������JLNxt��)��j�>eg�z�
o�"vO �f�!>:�'�^��mW9�o�R�ӪhhDd����2�.h�V\��U�S�ǁ�rG�Q؛�+{p�p�o�(=�WX�]ɧ��LF�u45\��HB^��OR�Tk���v>VLȫ�zbevD6{�D��i�VJq���G�(�� �$UTp455�Q�{±zfʴ��\&�sM�>=�||0]��o��O/_�,���"���Xnv[__Γ���c����e�j�ښ1"
J��L�K����� ���6-??1�$	i��͖�:h[�N�7����D�����n�e~U.@Y�CR �� m}��kd<j��s�Fķ���X1Xۢ*��u������_�FW�Ȼ�pr�ż�,�������f�$$�ư���-�R���j�rE�'|||���*י����!Q��Gg�����U��_�8�8� �J��7��p�,~P'rv���_{�]�/����L��Fp[�����������++�NL�GE���;opqu}�����*OUUS3,9� pG�0ç�j.a++������Htuu#��#d��?�aY���;99�/,���Y�����P��,�TS�O��S����:���@͋��V�)S�Ѽ�������-SQ=�:�p�:�F�}L���������-"����u��АN�ޱ'���)��Җ
}))�B����#��ɩ�N�77�_��>{� ��B��i/*��@.	:���E]}�� s���S�C��f<����ju��82	�������_�-͞qp8�=a#�����S	~�K����a.�C��_ �3��_߉�����j������������&&))y���JF�6�����ۏ'�p����BP`���?���'��6�\�����LME���ע�23���B�={@��񃪽��Vb �i�`��ܤ�;Q*g�SSS�0����;�w#�/� �g��U�B	������9b^�8�,��a���S{��S�R{��Tv�IS#@v�߾������t��v� �_�c�)sT����L�������!�1��V*�GضvvP���^)�8������C�n;�N�����t	� ẁ�q9ߒk����2J����B����=������)-�k9P�h�ᾣ�B�T�TNX&�DGr� z������'�ť9�!�ަcaA�0�q#ʊP�g�������{����~T���d^:;F����߼@���#*���(6 `U�ef���E��Fvus�A�"��9��^���`eeU�����Պi7�tE��Q~Y9�.����.`��d��񙚚B��D���*K�X����T��0џ�3e �N�#��DE��rNM�*� K�ғ�ξyoo�sd�{ 5<"�p� ��~�
>��=�����М���(���p��P�S�-Ԛ�hc�-�-�a�w��^=ssڿoC$���l >7j_�Va�ߥ�����@�[c1|��k��A����dd���	ֻ[T��?i�����&��`|�Qʞ; }K��T$$��[5Gs��ǉGr�l\)W� �7M"��D�����������1�A�zx`�@�w� �IThA��!PVٰ����:`�X��T��)���`�Wf��LA��a���,��U|���7�Z��,!�����[(YaX�
��QSs��W2_C�!�v���g��.7l��~������s���j{,P�t��E��*<���P��Z�1g��/���%��VV�	 UBG�����p=7h	��2' &�2���CA�q��WΟ�J2��"�mw9����
*�ꏧ��c�ߔ��3��-[��M�ϧ�v�3�A���=�����7�]�Ue��ˏ��:1l�y��2�����" p���I�;⎻s�;�AS���h{���`qEEx^mkk+���H�t\R�(����Wv�D��"ﱬ���[v�1�'�K8��춛�����(0���X}���.�؄�*]������x� �v�ZZ�xv�a����0�F�E�B.!I��R7}�IHw�ףsT�*&����O�X�Dr�@��� �O<�t�Vg�9V���������O��{�����+(@a`�Wekii���Ƶ�0g��/��Z2�~�����2
��2$H�h�ǜV����_-!��8A�[k v�|}��Y �X�>}���.D���H��F���oK���_x1�70k�&��OF���]hv+ҩ��Z��K�� -/���14��3�C�gO����m�z��wg4����v	I��*�k�G��;�]���k ��\t���S�N��R\������
�]�d''�Ǉ�	 �О�'��������[�à ��^e>��7q�m9�
�y/�J��]�����ԕ�1���l�wwg2솭$����p�hih^��,��Ti��ņ��6Cc~M�{��Q�9�9�z�$v(1���ſ=����R+�"̣�z��ɷ����?�]U�kz�4,�:�6a̹X���V�2�?hԑ:�Xm�B�qy�3��M�_�<�|+?\g�@'�ǲ����u���v��]-��ʓ�$�1�bT�N0z�ੜ��J�����`�������Xa�0)�;l�n>�3�m��.���9<��q�o������Z��z1���Ŷ��Sʳ�[���˨�7B��wx�O�л�z��7--,D�H��X,P��g�`�]H����p!(������G ��'+"a}��D�A		x0��ϱ�M����a�[I*� ���z:;a@�����<s>]�v�Â����	2'�d�@^���84�U������g��돵Âu�wszԸ��hjJ�I��վ�ۛ��?{o���X�������O���k�V�(��KT�!>5��e��2ς���`�o�C�L}����eV�O�-+z��A)��O�W�Z3_	���|���c�Ҝ�h������_UC��kb��va���\�OM�y~��׍ �~t��.r �j����V�'������Q�;�QV�%�p����#FGF���C�9�Gx}���� 	�w�WG�_�|���^&n<5�cf���� ���=�$U��5 �{".��YYY��m%��ħ�i�Ð�)"��7�m6~�i�������ٳguN��#܉T>>>���Vk٤"/$�a#�+I+��"47Dj�jh�3S�@$9���e��-�ң�����A9q��j2["����I}�!D�F%���T�ʊ�T�$<s�s�Tja� 6튵�L���m -sKJ�DDD�_�ZX E@Ƅ��6����˫D�<Z�)�v����V�E
�Q�� Ӵ�_�ɚxzxx����'�hށK^?��`	{Q�*��bM��$�"g�6ɡOZg��3KP���B�|�Z�|�F������^P�@L'nC�!�kq���K|��-x��m�s��U����L���"��;?�VV@�l�C�e���EDXp�{�T���S�aO,L�ys
@�?�ƀ�Eƺפ�˗�?���-�U��L��g~���G�ɕ��eǤ5�b�h։�֭���\����"�t�\F!+�]3B�<�h:��N����7��i��O�>ge-�͞ۆ���F��x�b���yՓ㿫��Ȉ�������J4I������g�f�V��b��H\s�Ͽ��nd��ݥ $d����or�'��@�$	Zjt���d("�T��݋�����t$�� 	YY�@<�rp�XXXx�^=�:Y�w�����*G�u��^7	z�@���r{ 9��+ ��VD75	$''Ӏ/@BB�~�y��{��TQ�A&�� l��Á� & �����/�|.,�nU8ԢR�����
�""��ZgpUCӠ%p�O�2k�i��"8����i�����5!���abp�'��t"�l���j��NO��8�hZ���r|��9�k�wu�x���@?�����49v�?a]U_�C��'���d����kp55��w*�� mq���9��Sߞ�6�tp��Ow���2���lìGff�M`���g��p����Π��ˮ�U��O!�&�@��tv落�!/-�9T��҄���	j�0:��K�?�2�c��"��/5�y�k'���l�@�WG��>�  ����{m�����<��i\f�߾=���+���r֑�w�O��j�!V�G��rsYVkO%2o.ww6�SYRb��6--�9%?	YOO�8	�#��7�Fc������._"��X2��nLᦖ���"��5�mw
JJ<\�γ���RVҞ��\�����[��spp iX{��Ԑ�kG� �m�X�q������
�y��������s���A^���iU���������o�M��Q�n�1;�M����??w�$�|e����D��Q���Ae�<O���L -�-������ޱn��*�4� ����"%��������J�7�p zY_2��Yv�#���m��~������s�����B�>ȴ��CT������q))G�&���������$�4㖶�n\�i��x;;�7��<�m~�оS��h�v[F��`MC�U��P���pQf�ms�l��㲲2h��q@@��J���%���f�/���������)~(\Aaz�?#�����?�검&�������CX3������6WE !���x5�^ ���?�6��xk����m:��@���`������ؘǬ�H:���i�_7��׷�=x ��r�6�ff��.�|����P����0��u [{ ֓p��Ar�&�W76�� �K|�u�v���jUc҃���"�ߵ�jD7����߰��捪�����@��13��qy���Q4p ��@K{{��GT����y;	�"B*�����Up#ͥb���ő�d��	~?��9y��׎�9��rOP�ݕj_1D�d$ͭȯ���:24d�s���8���"��Xl�e�I��֔��!?�gG�6%���O�̖Hx�q��?���5p������B�{A>;�BBd\\\Rb�M��#��L�В�a�ˢը��㴟�l_�����a���c�����t�{<)7r�t,��ȴ0�g�;�Q�� g��EACCß	����H�i��W3�����J�8
A:g&{��\pA�2=��2[��!�E�ET	d*�����!����P�K����G��#��Ճ�.BZZ6��	�-fff �����`'���$
��K�||ȝ�|s���s�teYĔ/={�O�c�6��0�!�|��/��*��s"[%����@h�GN.f�V��r��+�������..�(2�
X��} ���u��ݑ�����e�TB������͌� ?p��<�&|}���x������pk�W�p
/ٷ�F�;A��?�폘�H������`z�ݗ��@�J|�Ѡ��u$;�{�s	�ׯ_[��~h��U�щ�<x}?�������Y��A9���$-!/S$��vv�.9��R�s�O�<�AW::�H�>��]���Zl��7�onJ�X���Gr,\P�_�	�&��p+��Zr�34�n_ܧo�H�#�ǆ6p��]�����j�Cy�1�L��H��9x_iJW�bb9��]f�uM�88 X�.���O�oѓ��cG}��9E����˲xOO��9��u��x���@�+D����Ξ�JO��-�졣���o�_x��;�:�����n�"�to����9/77�������	˵�V;�N���\��cjrRjQ䋜�	�%����S���f�N��S�i%T�ӗ)�ʕ�a��49є	ޱ=~�Q���-(6��8H����q}�M�8[�7��sv�ү�i����o?xq�ӡ��L�33x��j�w��U�������j}ӃN��漀X��`���{��<���4��:dY%%h�O��c14A���ka������[��	�N�G�i�/F7R��`��\<�--E����`D*�Q��Mנ�S���8iii��!���V�ǔ
�T�9�x������! ����/t<<<5QQhK�k�3T��hlle�C��,��8b_>��@|ch�͚�rq�{i��I��OO�+4������j���'�����<�S@tV��_����כ�b����\�c�p����61o�B����c�����a��t2�\"�7}E�&y�H�ٹ�@W~f}��o_��_"���	�ou���:�ǿ� `a�l���9�ņ�n`|�ʯ-��hbb�Q�C��u|�&�2dc0*&fo�\�O ����P		c��&�7~��sn�������l�:�d���k�?��$;�x���~8���� #��^��:j�8���mm��V�<�vvv�g�>�>��~�j���z���`����L-�ͪ�XalVi����J��l�5	�yB9*pz�F7�۝�6�g7-Drઐ�2�AzI�eI���2���g�+$!�Օ<�	���t\쑇\0�������F��
'��3<��q�X���M�!�	 �Y7������0�q���䔔�dEa`f�>����a�����"%�_MU�]k"�]�J#�<3�7^NZr���V�&
+X=T�)E�[Z6�������YiKx�l#fhD�v,�lBEq.���a�,���w�G��h�����}}�==&&&��ֿZx�YR�|t |vu�k).+��P��1��%mpZ�S�M�����s�J��R4�O
�=0�q����ӝ��@�/!��-����Y� P������+��ꕃX@:ou$h\�>��B�A�.������b�0�>�pީ$����`�R��߿��=G�rm_����d%(]�"5���`	�U�KO��<�6ߔM���Bd �u��a�n-@�!Rw������㯦�t'~��N���w�T54
�')�`���ק&��=}��!�y�x))��� L�����"�L~��
�֐�CN��:��5 �㚸�nnЉ��vFFdj��g=ݵ��x�����;t��޾��!?222Pe�0�N��������>l��~����nle�/������?��߄ �zf���7��&�����}~~��L��Ќ�������UUUA�C��	��Q{{�¾"w����!����T"�?�u�p�����#[˸�֚-?����{� ۀ��ˣu��x����L ��^PP�:�jy��ʎ����o�;��F�T߼71��.[������Z3v����8��S����V(���'���Ņ�
��O�5�^�<|�0"{�A���c���!� ���[[�M8���g���h���t�,S>6#l.rVCY�-�C�U�K�PYl��nZ�2!ɿ�55�}��pim-�~#.^��������cNcATL��>(z<_M�M-:R�����`nYY4gy��c9b�����><�qk���C\S3E�@�q|��f|2�'L�4���"���z/��Ь,JE%���"��4�`v~iAR�R`2|��{��%A����B1D8�
��G	5Mڍ������8r����2j-�1$@T�z}�]\\�kC
�/��[�O���pf��$7�3�z��R=s�?�p�*��*����3�G9ĊJ�L�dc�e׃2�L�n�����x���l0m��ǭ�����toN�� �wdLL�t�z��Z�L�BEq���z�L����2N�����s0¿ĝ��a����\6�66ޗ��ȵ�}��u����u�靈�,����+k��I�,=��e�Y
��L@d����{�\.�2���y��
9-���@����=�5?��F6���ɓ'ЦB�7o��?��6q.��Q<�u��ٛ@ �h�אk�g���2�v��{/��T��&$�{�TU�����a��n��vF�3�F}�X䲼4�P�?���J��h^5�� �xv��&����s��No���|M]�]@���S�Х�P
.��0J-�d�c܀N�)���XAq1*����/�Z����300�
�z��Ѱ����<!N�F��7��J4X%$$ ]���(B�ؕ�p>�_-���²���9�^)\�̔kw3J��������O�{ވ�G�񶅻��c����V�P3�h�ba�?yrXD�nej�	p��M�����8_����y�B�>	���E�Ç�1N��& b��z"p"""P�@ʦ,K�����/�4Vʔ������3n�-Yo??�l���JJ�<��U򲼡�b�
���ިw�����W.l�XX����Z4��������s�����>$Ƃ�7����<��"�abXr���jH"��A���<�x��:�Z���-��M �n--���
��(Y��ȿ{�n˷�a�/��N�K�QZ�W��
�,�n����mrx-���C�6���V)�?S�x���s>��&�4~�L|dmP@�t����,�����j��d��ˋ���PUU}ec�Z���w�#0�N9#3����^�ܝ�˥����c���II�Y�Ȏ��X�_ժn=A��,a``�QQ�B���a���u������'{��#y&**�����~���c����bagfz���p�M��s^y9f{{;B�D�5
��֨��Ҁ���o��a�/(IHK��ov�e�'m�Afzz�����|��9�����(j:�1EΛ�
=8������~¬ͨ&t�ᖐ�<0'j�>�c��x���&��y����\��������\\
���'��?~ ��˶��~;'����E���f��P1�'���p�Z2����br����C\�Z�Yb���p�{�-jD��jL��������h��������l���SV@������C�Ğ�n2�v�<[m��uMR���P�T��CA˕�<=�~��<LI����#)ГL�YJ>!#���ɪ�ȸ���^���~�����ݽ����}w����� A�����߹��J�������<����3�� i�6uUU�����vR22�����G6��V�����'{{{#[����3�ă�n\�&&f���H:7�7���z���e�"�y(������/��#m��`�)((CƋnP�c��HZ�ݷ�]A�� �%���W;�?�A55|6���\f}�;�PO�R�2��("�{�j���݅���R���DS���������i�,#'�bW'�*d���T�������HILJ��v�EE?��%�Ń�ٵ>�ļ)+)隙I�u#�,N�pw��,�E�%� �����.�G	U��P�e/��x��a`b� ��G������x `n��QQi]�vFֽ)?2��[��]�6
��@N5���=6��X�7@�` �3����1��PWt���Uŧl�P��鲚 MlEy{���:fZde�*�if��J��q�>R#�������qh�)�J���~@?��2gyV���ɘ�iTRQ�sëUi������BmQ\����r�T�3���4�+���1���R22�g,db@�2`{���mtZ�1����"���N`�`���r� AQ�	��*f	���H�YB�d�������[HH�Ös�Z	���d(�Vn�����pA�B�BB��fo�*KK7��	#����vj��F�,6� Mr�J���;��O(0 ��4�9�D�mi��e
�����f������������0�rhz`�qS�c{�g�r�W0I��`D	}�@&��`{�h�|��V����O�Ku�� �ww-^'�5��g�.����y�X㡵9 sN//�jk��Ӽ�F�:��ϭ�w�*���˥(3���]pWZ<0���)�)kkk�ww#>��t��l�������!!B^ǘAUiI�%--dV�ٯ--����h88�A$o��Z��Ƞ0+_ؕ�}O5n4����� �Tꤧ���=7jgO��2�!!#���1絠�Dف��A�D�Z������lI%��	��0�@f
.~<(�:f���(z3`5P10��:RRR�n����@[���
�-�rXf����$ �J���ϟВ����˿?#@EQ��: 2P�Ѯ����t���:�a�EnG��7�::�@�2)e���H�W䆄��F�;"�_�~e�sc�%��g(�LK��t+v�P��hJ_�MhyxHʫi�Z�7����Іn�x��ʾ�EhNZ�������7W44A�6��<���z��[^Qwy0�	l?C��w/�Ո��������["v��̶���k��f>��t�w�+�M�?�0�X2Ə��@:��܃� ����=�x�;=u�*��}�2s4odq^=����su5�=�Bp0V��˗/��M�\M'�r22Н����3�ԋ�S"[S��Em�0�Eg�ɍ��|�dd�����C��?𙐾��<���B�$�4te�5�p"���2A*�߉*}s���?��*-�_�2X����u��i�I��ǌ���؛��7������C�S�BT�ZZI�*!O�9jB��7�ζ��KN	�Ӏ���t唔~�>Ӈq�0�d����f���@[���h���Y���K�;���80<�D�NZYXĚg������C~��$I��/��l�Z�K:��Y�0��)��}VAt
=M�C5�%� 5�FFG��lB�X�H��w��ɈAl_��>�� -6z����������ن��d�m���Ų��T;��=ɹ4a}p�Cj��0	?�f��,��<6L�Җ��L4�u�G3��!���:߶�'�_��0�Q�6faii��f.Bn�����.H��K!'	�s�ַ�
���D���h�	�6�9=��aO���[�|���V����46�WS�{�'&�X�\�'��\/A``a�l�rqa��_+�`�kq�����n>�/2��47#h�e`@���`�t�T+x�"� ��7%4}P��� �.1�`V�P��Å�#��j�mp�[z���L��,�> �I;��إ�n��%��yC�fڍtn�^�h�!^�߼����±o�~��wo().�U��?�QQ���	c�,�C&� ��,lS��
���͍�H����9K��N{ n��9L.x���JR�u��z��z���G�Rے��^�����@~A�hjB������)��Q�֡�?1��+��[롺&��T��������L'�HSS3��~������frJ
�.����m7P"O�ͦ��l�-68dv�8EEEAmm`�u�,pehƲ^F��(.-=��=8*U9??�ܽ�B)�r�%�爙��.ɝ����j�$	"2���>9###PDM�7���\����X�x��
J00�?6m���������J���@���&f*��++��UUC�CpkZ�Z���Ū	8r�H���oo,�m���?|������s`_L���7���U�%T�@/S3�)�o2�V����ID��}4�����
�'4<|�(����������������V+ˇ��v�QQh�߾A��0cs�9~I=ίi����?��?�Wc���l��T�l�%#��^�����ۏ>�込F�<UDG#���RUCCCo�1De@��:���Tt��*>�Ep�%T�oxx]W�Pa薏s��d��p##�+�8���˖iW��kx<"������O�Ww�#-U����h���1�@/̍���
F�&'��8.��F�Oޜ�g�P11;�+J�%tɻ�p�;�p�Y��dA���d����4�Jv�А��[ŕ�g��߇�������~^_�׮�����.���`h�q��Sd,9������~����j�s��O�"Lz�M~�x�6/{4hkht���Sq`��8p�����%H�<�e@'\`��j׬X�eI�Q<�ֱIJJ�̎�^���Gquu�܍���+u�ͷ��pӓ�6	���hf�Q�}���{b99��,{zs`J
N�?�� LC�W�	����x����`�r~���8AV�١�jp�'�����~�{qtJX3}̩�d4��M�s��(��p�3fʴk�e�ӸBx�M����fn>��Ή�^�,eEE���ֵ��X|���)�޾��m�N/�v ���[q�C�����/�����S���3'9�~�<2�n�� 1�\�6��{K�)�����uvsq<{�$�#�H��tb��89_ihd�	����8_�(U(��;�6�M$:��޷���:�]���g�~������-pȧT�Њ%Ժ��)�n	^��(YCg?_ck�/1  �	�/r�zZCqL@�? �W�қ|��or���x��?г���4�����������C�,��	� no�aN,M�(�k���3:������;>>~$��ݱ,�L7��;3 ���~�w4�V �O�q$++�	4H����kGU��I�x�ZV/������#�3*�� %�6��?���2B��Z�����5�Z��5evvV"���H����˰�v�l�x2Z��Z�j&]3s�F*}������er��H@Tɀ�! $�#%��
�i-T*H�[p�&����f`��~�t�
H4�7/�������tDf����0���d۟+�3M&���j���6^�;ť����"]h���Z.n�'6$�M�,y6���\���ߛ���c``\�ܘ
�it�l�_xϨ�j|w}�����V�m9������!���� ���8�ʢ���8;�VH|��)	�+�����y���p~(
v�`'Čo޼���/		����7ɣ	�v��y�R��S��HDNNUAm�pBfy�*C�VS�P��<0н/�~�tt� ��'� �j���>�������P���V�i)�>��W_�r9��ҏG�P)����j������X�uΌ��/��B���
���9a��	9n���#}v��Hv��ƳEz��h�L�:����5��jv���@� *�`\����PVHw�!@��H�,�@�(�O��r@k%��1--B*�2A$�1�;o�����Z�UP�!$n�ċ=����O|y-��.Ô�@2�Tr�Ҷ
B���h6����HZWm�;Bb;'zGG��G�M߉� ��|h��,p}�JҖ�����F2,�ar��ES�V���뚁�fec���[ˤ���`vo���Ct����4�q��5�r�b�kn^x�0�� e�g�~4�l�b����
�;�-Ə�Ǖ��z:\�ub5$�������CDA�J���ÅZ��[�oX�u�̟f�����J��5������O�H�%y!�WR���C���|��ŕ4K����P$�~U�_����Ѐ40�����AO	3TW��b`b��[]6��a��PQQ��������g�$T��u�"��M�����e�<X#����S�x{{Za��w1Qm&�/����kU]`"�)�w�h<H ��<�r�G���yaa
��5�/^@><���c�3 ��\�D(76L�1xȰ�u244<=?��wz����5:P:����i)O����Z�_߽LӉ�����3f�VV�~>Y�.�l�_z�I9�t���<S���bX�ύ���F�������J���L�,��(���T�*tz��8��ݏ���utt�m��$����}K�z �����QSScR��fq)(F�nANpܝ�SKe�32~9����j)��?����Y �Q����Mmچ�%r�3����,��@x���X�(x����ɩ>�[P����<ן�3
4>�v�V��Z����Ф㩰���!Ƒ!�������4� ����X�ht��ā��'$/�㍞:t� 1����0@@=v�4}u\V��6"!]ҥt(�!�}#�Hw��� --�]���t�4HK��<���_|�}Ξ=;�3׵;3� E���("x�����GIP�'ح��=o���}��>� T��(�T�	�U?�蚜��锾�)�;_:N��_���~�o��S�=Wt�7F};=u�?a0��-L���� ������-���@m H�J���ks�EXb�@)/�π/գk�Q�����X�>�y��5��4p�_z�[YI����<q��w�T�ݔ�D�5���I#���FFF�O�\>�4Ů`>��|�X=<�1��jV��~��)��~�Gn.����m ����$����>/f��w�����&��q� �8�N�`g7�� �{����=�K.1�{l y�N����C��|�&��;��Y�+tq�s2�[rr��b�{{{wu��-���p#�΢��B '����9 5O�m/,D �x�{��/mY-{�zb�h�������
����_j2~w���j�˱���&]���L����o`�
��{����H����d��W�@=><<�ӗo��'��G��J}��	��=�f��N�������//���S��j���wsv"���,z�q�hz|�S��`pbb \�z�M�H��E�ٶe�	�w���^ق���J���!F�?�g2�[�ãYj� m&pX�N�c�����������"&� ����HH���x��~̯|���#	�z9�
C�����_�7��2x<@��IIIu���^�Ù�4Q�H��ˁIKۛ�d����=%(���:�˅�-��i:7hI8�eý��(�(�����1�q6
��F]����<�߉�9L�U����}}y:󫪫{K��Շ�a���>@�;C8��I��!�Լ*BP��V�w��w�#���㋖����`��=�vGR� ���ޥ �D�W�'+��H��1Ʌ|wZl==y�Ix�cQJ��� ����,���Z��下L8a����lB�W��c��y��V!�7�!l�#	>}/�O�Xg�NƤU��$�*��=�_'~D�����V|�� ���q0�{v�ng(� ��,��2gE�����d� �öyd��Y���K������"
*V-�������@9$Mp�Wm1Csu��`%��jhb�i�/��t/8xx��RH9����`KW#b��^�����51�-��'@���N��qϻ�����V�)�G�t���P(T\J�M�3�U?�����XP^%hD�明���8}����m�����7:�JFcs�P�[ H���\p���$*u�!���&�n���t���t�3����<V:� �?��\�b�_H@H�����������װD E*����H�`�>>g����a[bai	��Y]U<�[&�v�����<bRS	���4����`4�,�M*�{c�0�-ֲ�n�0ٯa1�X^E�< �:^�DWUU%�|���7u���\_�\�������ӓ������Z�!n�بY
9�Ҵ��rXKL�� �gr~^2�Y�g^^���m^�
D� �f�_ ���lA�&)c���}D I�Y/b��:�#�����:1�-�_(?�4x|ږ�4�������,07���:��N��\�����v�����Elr2��\x82�6�/�<���D�@o��M �~���{2�$[7��`,0��y%�󝖋�D$��	��219�+*��Ec�LL ��l'p�D㍂�����7,S��+�Bx:Q'#�=?���oQQh-���SR ~�x̒u_�"����s4?2���E*�� ��o�(�D-.G��ٗ��#������B�I���0	� ���f�~�LIev�jP�"�����!��m��T56 �Z����$�q�����uk�{_�$ ڀ��m��a�� Z �襤*(��� ��� :����DaH/ݬ$���f��D
�����+<jjjRN�Q�� XX^�d`@���[h�#�����[YV������҆T�wD�����'�ݚ�N>>�T��� �P��Buu\ UUWwBK�M�>kk��T &4��O��H���`��kT��À���iEa���D��[������zo�6��ihs�JjV��
�ھ��Hn�j�ӹx� +��c�G��7kQ����}y�u���@&�[ڨ�ULw
�>x��#�C���ܼ<���vN 0P;����[[[�͜%�'l&9ykp=p�mt�Y�pg?��Y�t|�Υ�������6݀ԫ H,lu��I+�������~?���3 �Q ��_��~���l�����& E�
g(fL<Z����������� ,q�|�@����@n�f�`��䖔 ��r�t;>���qI�6oXހ�mzzd����2 A�6��住�������˿��?�|���T�E6ii{��+ |<{�n ��#����f�م~8��� �F�k�q����d� 2�Y$`�<�H��	>��h���P V���JŞ,��f���^"���S4)�F`�X�&�Z��C0�^��j��[0L�2��ю�Mv�[)���3-!2;��N��M����?�{��9<z���IO��4�����A�w�<�!��F�M�4�1xUs�P�8Z^���2�;�/�Q��GZ�X�M��L�����������lC�Ag��~�]��pސ���s�'<%���ο'g���20�Á���������F�I�j_�'��^i������MN��-Yn�G����?�-''G,�o�r'��mmh�Ԇ��6-Ɉ�k���cD�)�U��0r?,�P��[�%��v�ȏ�'y�y@����xxx Kk�h�F�����@��ڗ[�:�<%e�����[<�π2PJD
͕�&�5�D&�d������cJJ�@<�,�G�89F�ἂ,H�r8>��Z'u�ͭ�ﶫ-9N��`�%1��ٽ>(dx��\�gg�ʺo��7z��-�p�`���sB���%���x�cqi圩�pb����P(|�� 0�!""�@
�@�b�n�L�Ѫ��A�����A�!� ���t5(`uǔ�-�%�����Y�o�iO��H	�;/u���Db��s=�w �`�ziz�z�h��ę-vD�h�TvY��,I�DԤ�x�G���gƏ7ol�vh��sϩO.�����-�%z�G��o���ƹ

p��cf5��%e��X,��X'%�:�8�Q����Sڷ,��v4��\j�Ц0$�(��� 7?iuH�l�6�:�5�i�3�4��Ί�G��j�O��G,�����Ѣ�We�͈�6<�g�h,J�=	�6�i�̌��*N�H����"�#�4������&)�i��\^��1=�7',�yģ��g9�/�k��QHy�5A+�wC�=�>�խ-V��[�$�E��_%���a
�QSS�o���m�ۛP5=�<��vQ�٫�KJJB�"N�xr����!�C�=3����O���pW:23I�#bb�:E+�	[%$���fȘY2ϡ�/��CZl���Ėl7��Q����f�<��[�ju�u�ܖ ��q"K �t I���_�5W{{��~wԊL�:�3=0����q��
����C&U��&��#�`E���RFp�?`������/~�ߚS��꧃���Op}X��\�TfX/��󪬛�h�OK���6y߳�ȧ�)**֙O��E���ۦ03���8큩�緷�t������.�l�!�S��,�6\��B�]��Zq�U��n�ݏ���n0�K��0�[�	�@�6Z�����5�����N4Q6�>�P�x�Vד�P,J��:�`~'<YY�2����W�_5��}k����u�L�u-,��V��=9���n��U�@X6�u�E[����3�r=��D�Amw`�L�5�P��RË���@���ΑQQ`0\$�L��vu�����zW���b,~sztv�!/ۿ>III�c���۫�*��ܙ�"�<������[ޡNMM�11հz�eֱ��l<�UvF<sM���f\.K#�o�F.-��P�dĵ���MN���(VD��pMůj"}}x����� KjnU�P�Ϟh���nR�WV��8�����p����l�>r�m�^C�T�I����t7T�=b0DZ�'���PC]���� uY0�`V�]��d�J����#��t�.)��߭i�F0���b�~=~e��G�X*|\�&&��xV{o�)���o����4�yAF]�d���CC���$JA��6��jH�s�N���Xd�$?���=��1�9)�	���%�$�ֵ�`�W��+'���zB��|Ê�w���g�pREM[�Uq�p�O�m| 8��t�y��-��ԯ���y���I�T1�ϩ��}�)(��wv=L�t�~o�7	g���=P�
�S���7��01a\\Nt������c��	 ��yE'�?����(A ������\Ȱ�V��U���e��+<b'�;8�'0�%u�*���h��K�EWGߐ�E~]$Z�9�:E��K �у���( <I���mm��+�p�8������*�A�`� �:8�ZZXl�u�H ���G�Fr~�w�>w�K'�?�;�[X�/���t���o�Q�����ܥ���U�[E��w7eML�h��"����|i��`�z�Pcԇ�x5���>'9R�%�/�-�K��eG�M@OO�����Z�wor
ob�<�Ծ�&��P���K�0T�����ɉ2ʄ8W(�
�Y]-8�u����ͼ�?�V�6��Lu*k��K:������.u�_h(����z��L�$���Ó�x{�> f�,�uvMNb��	U�=ܐ�?�V����U�D��J"E���ӈ�I���/�:�%0�ދo4������cŗ��۞��� 1�/(����B�x��947��X��~���T�(ݕ�p��}� ۳ ���$\4���gj����A�Jb	'�"�@��+i�g��d���6r��_�fvv{���OH���q��(*/)
�[v�_�X�k_�!K+���w?������0�FV�n��6�y7�.�iaVF�ERE-1�܅vA�������{8}��=r1%%�:$����\t�s��p䪓���f� ���ޏ�y��ƗdD=\G�>������̙9�^Ȧ2͊�H� ��K�8%@N�7g���d�_==���t��f�}�z�}�s=01���-"��O�����xʱu��u�s�J�!l��9<�r��ү�r�t!,���,W�'="��2��!�S̠�Y��w��n�q鷧#��
������!�UŭPh7�on��6���yj5Tz�����_3�(L�.�Q���}F��Ԩ���P���_����K�M����#Q�ق��?>5y^3��`EP�T��^�o@~@����7�f�5!�V�Aۭh���e�*��wǾ��n�'��� ��\�tU�;{�eyu$Q���S��+t?҅0�ڽ��ٷ�����Z[�ՕsbRR���kDt�8��� >����ņ�l�ѱ1�o>=܂{Z���U�� `N�]NBM������*
�	���p��9�����2w�Pى����|�d�{}s)�'|��Js ����o��S����qx���@o�u�jcpg�V1,w���	n}y{{����Z�zyXYY��m��F~�%��3⩜�j�\���H���:f���`vv����^��¢ҡ*u;��!�K�4�M��ܨ��w�v'��lG䓛22��j��?���%H���B�����W����H`(C��69 ���N��Ů�4�p|�1T��aZ����=�IXS ;8���p���A��� *-����Σw	�g�������x���$%O��U�ƞu� �t��EL\UWA��C�Qv0�a��i�0�R^�*T���|�t��p��#��_|����ɐր��6����f�*7Z��!���W$ٯ�nj��=
�q@���/b�;�O�P"##�445���)�	��e~�4��0K��
�������ˎ�]�
;����n�M��^��
���u���%f������!�'�m����	҉�5�?+>;�\��ʓ���b�s"�d�ڙh�z"3j��K��=
FK���Dy��Ʃ�p?k��x����f�G?�X22$����㯨/����9Z�-���$�f'�e����X��j�px1c�ъ���B�"�ʨԐ�iܩ;7��Ņ�t��Q-�
ӡ;19,*�z�j���3X���'ˍK��|�((��S���"zΞ�������գ}h���Ԗ���a@X����E���u6�����������F~�{:�X�$%��}��S7�������k�����c��<C	�N:/�A(���=���ji�p��gS��/'e�X0"��� �u����1�{o���R3뵅��60����OK_k�2X���Mp\֔y%�3�|�[���^�5�,��A�%∭͑)�X|��=�]O�E_���ў�(l��ܹ��9?SL������0�����tL��0�\��L�5m?|�Pe2���v�7�(
�Y���1q���᭠򫩩������a ��=�����("0:Y��(��{�(FBC��\�0(��0<��h����p��q� 3w8���:��1q��`Q ���
���!F��&069����(Ɯl�)#'��uWZ�T���������FB�Hُ��-����ߟmʉ����1�SL�%;�3Ruw�s��X�ȵ"���M��K捿��r���w����\)Ӆ\��o��ïbù��|W��^6�쪰��=�<ZV������\,z���:'�Y� r����a)��� �M�|�p#��<�������#r��i�5h|�0��c��,K�Y��U:�% �\���M��࿌�	�QS���*7j����������LM�Mg�Be������O4 ���%EdTʗVF ko�$�UC|#@F�pLN��M�=O�y�p�d=���ڜ�+.��E.� �W}�%&x;�o�+�pc�6�)�T�D-��ncx�f�����-��c�K������^�b֩�)Z���I��❐�������Jޫ�(�y���Z=x���i6#ڟm%dho�|��,��+�!74LŔWVJ�ˣ����fgǠ�3��5��lG�p���y���RT߅�	���VQU�8(�޺�?sMς���l��8������0ē'���ڄ��c�����������}��߳����HZZ���b+�����*�duu� :�����M&N
��* ��Y�而u����PVFXI	��mzf��b�kb�4t޵��,Z^��>rHϷ�F�¾@a]��½��	 L��d�(%����� ����%�IN�6�	�|��+X��1����6S�`��hr!�v=�����	�\�� Vuy�9i%�V6s�qp�}�M��,��`~e���\�gd�����>�1�<�UWca����߃�-'�?j��|��#&p	�> �Gx�)V�𪅅E���Ǖ��Ф=7�]�����{:�R��I��l@^���,�lDyX`�-@����q�� o�&��	��� �7<<l�@�˗7\^��{��2�:��[����_V�Ӗkk�����D`e�큘�3���SPP�:�Z����w�2uKKK����
���VBUG���iM���~�� ��ć�_}+Aɴe��dxbh�2�Za������	?tDDD��V��j�*�g��ƹ!�@q��P�_�υ`�P�Ia�<��{"8_��'i�u�f{;���e��?pMD-����vܶF�}��Xo5�$�&]`����)z���y���eϞ�>����k�V��Q��=��)1K�����]y\�v[���W/�6�B��4�.�$r�����x�b�zsc�Q�ak�^�D0�\���YX�rr��x���7:K�W�n�7=w�#��{��q}��6i� H�r��#p����2}a��������[s��0��Cp��g�Uɐ�i���ce�r��h'
6F��ʲ�>ȥmD���R�	 g ���(dH�/���*\���˾�cKx�P����$�	�nѧ�n����hyS���8ZG�d(X��nV>���J���oM^��4:ޣiS0�cN���l@"%(}���K1� 	�U�=��J���{ׇ?	- ������/��A-�7����ˁ�}ʵSL��P��㱷��J�FH�6d��������5�{|����$	�����i��G��$ ����D{�1P��=����4z���kT�&ğ�e���јhrdT<<���S}}����3�Ᏻn�lk�I���xH&�v2Ix���Ő���r���t�b�ט/�f݁HfG.�ҡ�Ā�GP2�F����u�'��������lR��1�SU�&@�/���"�52���Lת��m�x)�}5T�/��#A0gm-.0��ƗإmuB�'�����Z��{}��|����R�ru�/0��!���cϥ=��u��ݯ/��"�T߿�g��+��~�۰_V	�O���	��T�B�J�F!��f�O_��[q��[{�v@�[<Pm�aL<��+{/u��p֞7����cSEP��5�,�,�X�V.ώ�љ'��=��	��7�G1�b/S`#�S%��h���-�g�E�9��7D6�\�~���Y���R��2a��-^���gX�]Y�,�nD�_@D� �y-/!��_M�y���s��� �e
 �m�ʟ?~����8��9�=~���;������Yy�nDr�s�S
?;i�|,
���0��kRctC��2v��}I���E!8�o+�F�!]���}�U��g��37Ov��F�ҽ�gbnd�T����+7-�ApbzF��j[T���^��"\lh�$%;�Iid2.����� ����J��0J���P�S����gec�B29��,��>�N7u2�f�]�;>E�`jWǏ����?�R�x�-��Y?��r���<9���J�s߰�o�/�b���}��o��`��
���z�pq͵��ܡѿ�$���	��_��\a�~ژ���n�Q��A�=-��Sဃ��4�T�:Ҷh��Z~bnʞ��?=��#91'`g�$C�/�ጸW�ǿ�!�<BO_K�?g��hPv�*�ˀg?��������q�L���Bi��	SO_ZQqsjk��7�8>.b�	��n���J;r�������&N�us��R��g��v�KJ�>jVώ�q+	���_�N��&��#��mi����}>��e�3~�˿����Nĵb	����h�':8�;������+���
�y��3=H�ao��l��	6��e�7��rnX�ho�V�{�����>	T[=8�ۇ�l��W�ױN�T������ͳ���%���ڳ�n��ڵWR2�F��\Fm%	�(�1��G<���:_sN��껇���=��a�a�����v,Უ�!f	�J~��m4$�Opw��� l�����Xx���L5�倛�3붜Q��(B�<����p�L^]�0�&��B��됕=��ECj���������u퐷�x���T���1���� :vp���o` �.�2���Ͻh�1�ٗ�P�&����c\n���jc&��g�g~/��׼����8F?D693�(�W[�Q�Rl�s�
]\w0�̋޳t�H�M,OLşM^�v�T�,$3i�����F���k:�.a"��no�-��pb���fG�2�*�� �/�Wv�𓹲ǅ���oy��\���y&J���{��+��O���I��l��U�n�ԥ)5�k���{,���HL��--9�1Fg~��sr��f��Chi�Crc��b����[j�ݒψ�VP�j�(-j՘�v:su����3��D	t�A���� ��!���/�ήr���J)�ht�f�;���V�k�=�������Tr��|���q��=S���n=�h&��?���S�x�&e����}���N�k�(6��U�<�q�P�J��`�1�::�4�(���65�S�^o�na+*�����]w��Z�$4��N=���ʆ54]#X��zta��Ͳ��ɧ��sN^��A�4�����yܱ�|�(��Ak��0:qh��1V���L_�)�5gm��Q̾� ���<�z셋1
��ڼH�0��$6e=͘��J.N.�/�?̗�[�Z^��\��$��*D�fQk	4[�3!��k�qIZ�6�� ��\��d������;Gֹ̚�^��˛���l{dfI{N�B�i����^��X���1сi����IYyр-���b���=?g\ֳ5T�2'�D�w��5���"�� V i}l0Xn�f0B��qNP�E��O�dwu{+)-=T����{���t���b��'�����Sb��;A����3��Rc�P��|P��bp0v2{�6�7����` �������B�q]�̗�Kb|��ċ�6"y:�y�d��L;��S7����OXXX�0�C�n\!h�e����ʔ���Q��G�!�����Sr���� �?Qq�憛�կ,��6_��>3�'�;9,`b���D���=^T
}V5~��+����
>�U2��/�$�6��ċYw� Z���[�ǿB2���!ɽ KW����u�I&&o�fJ|`��0���Ў����t�5��΋YON�������c��K$�ދǥ����|�Fxx/�d�P�;�덺���������S�S�j��{DD��sl���� 1�R��z�����Vr1QF����W�6�ߪ�}c8"��+��~	��,8���m|rpP�F�ތ�"����q$t)��k�8�G��SU�ܽ	S�Q�����m]���4\�O��&�ۏZ����bmO�I>��� ���4����b�����0�4R��G�}K�79�ǊZ�)�s|/7�K��v�!�3���i��Y̴2����`ƘHm�q�C���7���{y��SQfɽ�4��2_|�?����+s�����7/ՂW�En�z$�mm=&�����Ƶ��Oԫ\ok��WA�D����a�����S426�g5���)!���I�H�̡kSa���1���kcK��B�X@O<Q�Tԁ?�Lk;�����al�x�J��=��ωz��F�Z��G�7Skkҋ� 徻���d��0@x�d��XJ�����5�=�Մ�g*��[�ҿ𢐙��3��/R��s�Lkϗ�������U*�V_���ɨ*+C�sŗ/b5j��jFFfLuCU���ʵ�����&�4cB���=ZU�����œ
74�[�6�Z��Nk�g�u%��zx�@��\�Ӵy���̸(7�)�y�=�m��T�&^�-�*���e'�qq~2�.Ǜ���]8���Q�O��v�1�ta6�Mp!f|�Ј0��=v�~��9��S�Հ\lyͤ_����r��"�ܥ�\[�t���a�>jq�7lfb�W6V@>8��ޞ��&��_����s�Y�#�g��e0
>3��#*8o��ULc�϶LO�?��8��M������Kegt�)N�+ #�������_sm� ��x�6wy�3���;,�&�4��i2x�W���8�`�'5f}�$�S\�w���<q��L]�0T�)��VnE�9i�e��P%���c9�w����%M���E�1��[tN�쬳v��-�9�kBՏl%���L�?��g�Mv���o׆�k���06�Df���*	��jB�[v-����6���!'�-.�R��.�J�-�uPV�^�B�W�V�(<|׮�%C�}�
�{N^k=������l����{Ƌ�^�g�	t��M�<<��E�k�ޏ�2��cu����A`�������~�Zx�-o��`��+i$����F�T�ɳq�O#?�Ykv�O�I@��,�Q7ܝcDjN��I��јnt�3�W-�W���n'�m�u�� �|�-F��ߜ�=[��zIŪ��C���Ndiv�����o���U�B������+����<�_����T��-��1�l��Ƒ5�+�6�/� �1F��du��__���*�g�}o��2���A�$�Y^?jʰ���1g7ǔ�(T�/и�xH���ժL�徸ʸ'A�Ԅ
.��>y� ��>����?��V)�.9.�c$�8?=(F���px�؈nr2Զ�Q����QC�������a�I]�}��]�Rr����ل�:>m��G
����j�+�tM���?�S+���n	y���̺�d��J��A�ܽy�Q�^��D  pB�=5S�s%�ϩ-�_l]<~�(�K�=����A����S��8a{;4K�D�5+#Ht��qr��&���D�j����e�81:'W�Ȩ/�81����S)w^M��=�%e��tbgc��ԦHm�Y�^sVP���Q���"L�а9�7�Ez�w0���=�%���s��x|���2vbב���1.�&F�Ń�PQ�WY`&�Ĕ���X\6������~T�Ĩ>7�F���W�W�yE؈�h��`���nȩoQQ�v�Z�U"^��E�� ���e^{��;ۧ����J�$FZRI-���� �Ϣա��鞰N���rp��ڤ���7p��K��H�����5��%7ye�"�� ��bs�@׾|�ET:c3d\����!����� ���B=`���mx�ǖ���vi��d�vK���<w����Y�N.U�s}�d.�向,�%����DOں:�(.�K���gF+�Yq������'�j�ec�2''�w
8N.Ւ�6����n��_�.��פ��N����5TKtU��&�U���_'�v�`Fg�6^�%UR_�d4Ut��.>:�X���f�[�D�/+z(�t�k؊D���qh_�F����A��eq��I�<��A��N�����:��m|,�I�3
�2�i�x��z�>��!YV:����8��Qy^�E�ˇ"��_���\�7��망-��Z��d!Z��#���,oߠ;4e�d�`O��g*�@���p��S��f���T��J8>7� V�0)ϫL��@��O���%�H�T�����qq�����GR�"Ux��ϭ.�q��}|ښ&���>-f�#\�:��&��>7�����IQ�sS�kz�3'T��u�ח��]���}#�s ��Ҍ9��p�KC�m��M�?aˏ�;T�l���gjyb'\f==O^�ȌX�ឰ���63)�����YU��h�$�22�����4[WRnw� ��p��햜<�Rr��0Sg���;��0�|���;�����7���7\e<�"��ai��bK����r�!3�ң���lp��2����xT*��/�~��#k���f�j��iyݰ�3����lehI]]!��uҗMִ�eN���,��͔|�QF���c�>Vô4���P!���]�!���8��I��թv*��h���ISy�͉��h�s�222��cFvsk��x��خw1��^��-2��{EPU*�u"�����m�ȯ����?���b�T�k\��7�V��K>�'�Bu��Y��d�{n
xZ�� ��:���:e5_�wwѓbᱟ�VFT�:qU��yz(���PQpt\�� D�y�x�'�w�/��#t��!�%Mf��ך�NU��-�D�-�=5�����Ȏ{]le��
`���M��5R+�N�����L��ʒ?��|�����l��Д��2P���jib�/�r,go4�V�h��=��V�L�ϑb�lO2f��J��h�3��5_liZN#��5�k��WX�!�j��A���i�N-���R�r1|�T!L��"{�.-���Ι�:ڒj�i/	����*�ʞ��;����Ua�4[�A��x�eΒ4�&�GCy�)6��3nw�g�[�I��N#���~{�0Jl�K��f8\�Е���]��m�y,m�f8��G�O� *M�oܩë6У*0@p��]Ne�7P�B�ƓLe+n��L��o���5�%��&�r"��KmE}�l��-A���2sq�����XV�<C�r<ly�͂
�O����L<g�a�1��f���t<I�_���T0�'���mPپ�y(f�K����%iː$�n�0�h��:=%rfFȖ�3g���佨��pyϜI���q����M�R�E j1��Kl��FKfx=^A(�@���]3��kV�{`ϦA�ʑn�,~�ҒӇ���X�W�6*b1Ym���in�i�ﾏ���C��U����*J�8�^���EL�)fH7y����y�ZN7�0'�F��Ū�BD
T�n��|o[?-��9�?}��%�����v�ɯ/����r7 ���!,��|��q����p1�J��s��ںb�;Y��&���Yz���S�+����w"%��&���ּ���ww7g�U��挚tГ?��'��X_Jpܷ�M:Zt��L�!mj9��<cM����5.ᰣ�aƏ�W�!��^��L�`���z����؛J9
^���F�+U7�7K��TV؜*�2f9�@\Y�i:�7�{wZ{YޝV��`nyL�@���3�I�NvF�ާ�i7ƽw Zs����Br��*f�,8�������VX(�_@�H�En_�Mszog�G���PKYW���덳R/�8���م�%"�r` �v�y\�CS�32�~3��������G\�6cɡ��&��:�Yщ��vn&�(o���4Ä�n��ϯ�2�E�;�j�ҳ4�:o�23e�LO^�q�x��9ds�(z��9#�"��,U�B]�CWұ�������Y�?ϏG(Sń}��a���6���-������U&���2�yˎ�E�Yr#h|!t��1s�
��ce�~p1F�{[h�Xi)��ȼb"�Z�?g�g��Ո|�;(�"!��W3�w`"�����m�j�)*�p��v032S��@������8�����\�2M���ɶ`wjZ����0ԩ�88JO��K���6�c�*�H�/e���~��G�8�JKI��޿�����!~k��q$Zl����W�Ӓ��EPIIp�eg]]k��'3���/iF��DF5!��B���c���/�/"�6�9v��Ŧ��~L��Сm%[_Z
^
L=�_/��;~�;���j�[[�Ե�r�7J��We���`5��n��K����~�@'k����f)P��������J�n�|0��b��� ���W���\C�K����il�A�����ٙ��ۺ���Ӛ�*�$��Z��Ԩ�˅%B6+����RvC�4����T435��4ι,έ�v-q������ZxǞKc"�r[(_��Ffs1�6�Uy�+����tn�q�ʍj{�&$�m �d�XL� �'���@e�N���G�G��Г�h���ޕ ���35ޱ�~Mmj8x��p�1��urKE��Ăweɕ�D+lG>�kؙ��d��u��Pc+[��R�����X>����&J���ҟ���Ӛ$O��r��ƒzo\���+�I�w�0��
_�s���I�������]��4Qq���{�vi��VQ��0�����Qk��U��p����c��no˺XM��#7�Zۢ�`�d�~�℀0ʆtm^��xG3*����
M��{Mփ�a���bY������7�{�䢐�G/�Z۞ɷ���Z/Y1�eg3��#+3���@���fQ��K���Y�2���s�&�e��$=o�=`�_��kPNS 9ѧcZ�Jb�%Ol[�ޕ�Q���ڔ���#y��E8Cw@��$"0�~V�R6i{UP���翝ԛ�ݹ/#h��GB>�`���8�{<���B�����G��z���ΎђU⊂l�5��#�(��"��׻���?1��S1+��.�����HH�*wY�D韜\Vfm���82tuX��b�T�Xk��g�	�(��Vhӧ�Թ2�1$�*�8J'�qs�ϓ�#^�o�&�l�jb�1��|*t{u�kUَ ��(����N�pR��T٪�;)���BM��N(C����$0�z��C��z�C�у!ԛ�au�77�-:`kأ�$0VuG���AR�э����|6=P�M�s�BH�Mlr࡞�����o=��ޜ[b�[������nwU�nu���&�`�i��""4�Z����+/m��ܜ>�~F;��/jű<\(��L�)�{isf
�FNf�ۭ��i�=\�%�Pz�Ծqz�ϋg��P�S]Fks e�m���O�*��T9:��s�������a����s��.+�����K���W���
��RSs�j_���ywO�\�8`C�����]�ӡ���0HH���&��+Yß��]�"�w����I�謵�����c���f+6OJӻ��"�	�T�|X�Ng����9s�Y.����n�`x�4��g4]B�%u5��Gzj�2�!��7Z�k+JK�|���e<�^d��de�{��'�49z�7UĦ��(�a��1[ƙiF	�&MX�s�^/�H"�x���]B�]<).L� ��@�`���Ny�:_�]2Je8���_1���;��Zē�b��Q� ��]S�4{�V��r>����R���m��ˀu|�DB���ͣ?������}:Y���>�Ih �e`d�;[��*:w��x$�)����Y"^���e�Y264�ylP���Ӥw�8v�,��o�\��V`�Q����L��q��^�0;�P78D5f%w�U���yN^!�� ��|Z�;Z�D����B�&�ˎ�-L7�nr�W�2I���b|TB������}����<�_oucqtt� ���V"W���\�٘�"8���8�J���9��z������*p-y�U�.��?zz,�4��F]�՚n�C��&��<A�zY�� m�>�#4X��j`p� H �8C���ÿ�'�zF�Y	HH'n��aV��������o ��y½I6Ɇ�ٍmsc�ƶm�bgc۶m۶m���_�W��Tݙ�QO���9gzg<s�/��O/�;J>�z�q'���|�3$��R}�B�B�V9�SR�m ��m����䴃�1�~�Bk�!''�?����e���{$��	���83�!'��lx��l� 4E��@FUa�c���Ig:���x�J��A-�}6NY���
3*����B�ew�(�b�p��2���G�Y����%y :6>`������l���d��*Y�Ȼ��j�� U�v��L�M��x���o�2�t�i�e�0k�8��I�cɜĦ�%��$~��]��
Ƶ����d�A�a6DOxH���/N.���	��CZSV��;$nbpX2�&��&�.�)ٚ��*�h�jB�S_��=��6>AM]]g��D�ظԨ,2$u��SSy8��:޶���o�Ƽ���?9�s*�<�̵IEc٢A!Tf $���G� ��Q"��
k7�$�a�!�6oM�6{*qo[��ֱt����Gu���dQ�ݛ���YK(��&�/A�8Q8X�&d �А�>g<�J��t����<2������H� �U]2��kʎb�P�+lq`#���&+;^(�^�s��.7��|1���+�:�th���|�}7h��Yh���/��`Op6�4���{l���k[% �!F{]mq�$�tx�Ȃ�F�A �$߾<�OKP+�y��|����K�k�<	0"�V�8�Z�̊����L�w>���Hc5����m����*�Bv�����������0��"�h���g���gE�WH@%
�[?!mk�L�s'�NR�ہ�hP#�Xx{RkT�yu���!J����x2x�0� 2�>)K�3�u�3R�֗��@`�,ˡR�Lj�\������6!��w}���� �TJ��)�Կ�a0qo��H��* ��j��ܼ`b�@d�7ffV�Ѱ{�C�͙Rd����� �$u�ꊣ�Z5G��IC&9��;�� �	a~�����ǒG'�{+V�p\�|gW;H�u��!2H�T���15�� �d _�}�T���'��|�T�'t%�E�{Z-t�����K6��+�q��q\�{M5d�AB;@F5�F��e��'�� ��/���WI9� �x�M�Z��x{݄]up��
����2sc�d��8�y��I�V�rm(�s5������f�D�Q���#���Oc`���[�Q<8N��Z��j�U�f�W� DlN���F��Ոb	�)֠�� HY��Y���?
bj�r�/xʇ��P�Y*O@�,2CO�h�.!nɑQ�]���Ak~�ٙ�3�)4�;�V�xET!݀�b��b���c�Ydɔ�9��T�-B�G�))��:���ݬ���ܴ�I0	 Q��f�L�����3�b�@�iC�̤��T[�X��4&�,[$�u	�!Vr�(.	N����(-�������Z���z!�yA_�	ʞΰ�����m7S�_�Y�UMT�r�y�%ye�s�L9Ʊ�}�Fhh������]��Y�y�93T�_������K(f�D�R�KfRnv����ﬅ(>��v�����������}�����k='M���"�ʈ��8e�����{3��?�s�"��E�䊅�f�s܃�5:ҀZ*e�D��P;����q�s����K�i�Wl>��i�2�/��pA��{�2z��<�Ef]��>Ӣ�]y�ۼ�'����+��e��ߌ�:�fgo?�ml�S؟ݛ�4�)�~w�8c@>]�J���;κ)���:/�WW� b��uʡ��T{_�����Be��G���9jN�[��oȨ*�C�ĺ��;�7!������G�k���o���#�(��l�D(g̫��2�K�F(qy�L�!�|)�yU��ɤaB���c�߳�HKpCHP����:.�)I�tw��՗��s�g�$��[ �W-�o�=�&MާWc� �QIAq�:�e&5�+6��9R�B�Xz3�3�RTn�k%����tB�ԥ��U	��bs"�����5�)y4-C^
J\�s"U���a��"����3T��cGl)�0%���ݾ�S˂�no/Ɉ�J�*)I_+d�U�㶒3��f=K�[�?�/uz+)< J��)q��M�Ԃŧ]]��e��nſ�2AnXJJğ]�υOHA���d*H���,AL���5�@��$�b'G��ye�~щ��oH��2W�F�0�F�Aߞܞ$��m��7+�=��7������+4���'	%��zs-�CV5����pqV��I���^y?�>�ҍ����mģI��bv~�$�g���1?M	�viAe�nĒ�q�<o�5Z��/4��^�|���v�i�t��5���''�p�����P&����My
��ǕK�������;��b84՟�����:<���2�rgN��Ob�w.SPm�V(�:7 Q�k��;�'��cο�&��y��g����ߖ|����'��!�����
gA�6�����L���N��4b��)E��Ў��ޙ:��k~��� >:b���1u>tp�g<���b���65����D�E���.i^��V5
Y�Mpe�"w�Z������Vo2dy��L���1k�;*��Ɂ��|3Z�4�@��"G2��\X?���%>�D����}{��A��>|ơ�X��x����-���&P��-9.��'�&��?�
m �%`��0����|{x�O�F�k{���Ǝ��MCf�?�y��C�k=�,�78��K���gw���۾u�}��.�j���R���������Z�6�`|�b�J���;)����U����6W�쎷$`i�$O؆�GQ��F���\�Y��ށ):\��e��ʷt���@M�/�9�<3��A�\p\�(�8?����m���ɑ�f���S�0a�b`>����f��K}=H�eϳ���@!��k�l|Ki)�Nr�������_�1JĠ3.TY�u��&~?�թ%�׀�s�D��~~M%�[?���_X'�+�n�U�xh�]���s�ל8sHB�%$,�N	�U�4A�	��
�CA�].T�Y�:W4�� �{��w*�#Ȟ�"\�Q��k��tHM��q$��O,,N~�R��z#��BJ��vyq!k�f_^^^(`��a���/&K�/m]er]���H���c��C��3'�y�9�h�y�é�,��h�^�[��GS|᱄y`��c	�.dM�P4
��H-���G1�xV��9�"\�%�QY�w w�\�93C��������퍯P(�w<�&Y��s�\�R�V���f�ɕ"�͵I�?�:.Bڏ� ��Y%���O����)�;�G777�&���Q�諦�v�؉�l�6�)�Zx6�	
��V���\�vYtM�4�͓�����2�煌��b�j=��y�B3�N����D�U���8R7Og@����L���T��E�����37�v�7Q���X�m٨�R�/''f�+��rW�V�d��5���gV0V��>0r<����>ҽ�Γ3+�-3�4ѡ6 �P��e��Xc�/魦~:�T` ��e���A�0�_S�[T���h-��P#��mh���)����5:F^v d}Sǭj`I����n��Ɖ�ssRt������pw��y��j��ײ\�nS�98[�A醻8�I��"���qSf����Τc��K�;���r�D8��[V����j���p��6�fKC�Zf�Og��RpZ��m����7��orޏ�ܨ�t��c���*� �'S'��kxc8�
�:A&�!Vuj��bV,���Y]��b��,���jtlY�� ��y��� �t��M���./ǅ�22���W�gw�|!\@|�RD#U��1hgz��7��,������vH*.�0]�=�ii�q��H�����c$���vX���MȎ�J�W�Rժ��gC(`��� 7�m �;��ٓH(Q�;��.Y�Ƀ=�^(�[�Oh�/[5ؠ�_�G�XY�&�5XG}����poA~e����\�ޞ��vĄ	��U�Ab��Yp�#cC�ũS�߄�i������l���������?%?�x+UN�g���B�]�z`Ìs�)R��؉�w�xM��'Zq:P���=���EAQ��,��犉0L$ԝ�/��0#q���"R�zha��X2�8�\�3�Ռ���0��`6��	9@�U[F~ �c����c�Q���5�Ә��ί��	�1�K����wQ�0h�� bp��� �L����OP/�d��q�񺃑�lGSU����aR�,��V`��|��=
Q�F��C�|���<w{�CYY?���`X��puuuُW^����s���L�����v�����E#����*�ا���.��z߆M��瀯e!g� �I��<���$	��;�Q�ȗ����<=� s]<V�����i�6�g�'{�����G�)n��{��N���^5P����O��Ԫmb>��<Ֆ}9��yj0tDJ	ʽR�= e4��x�r^�㔾>��"<��,�(:��<��g(�|D���)y��+�����3a�k���k�E��
�G*?oUi�F6�?T��ٻvԭ�h��Xu�P:@ٛ���,%V~nW�����Į��A<B{�M��,B��/N�Yq���u�=A3B�L��O��mKK!��r�*-OX]� A~��z��E�F�N(��j�}�"�.N}��ޠ���OϾL�&d��� �{7���Vx�n��U!���ǿ��yxx�����
��χ<](��a�-?Û�@��"������=?�]s�uO��U-�l,� �޾�!�ScmU]��aT�б���&ņ��c�6��'�*r}��i��b����f�bf��!��9�W�O�|ۥ��	jf�d9�<=d9g���`bP��p� +�NG����z�ʖV�h��@Q��2���g)R�b��$匽h���~T@���ؗ*RN�:"���BiI�H9����z9��x��(�/���P�v#���*/�(?�ѳ2�E<#��E����3�''bb��V%�����j;�9�נ9��IG;����e�0�ժ�@���+��@�?��Z���#O�����̗(�+��p~8[~��ܝ�D%^<`���y΋~�:Ȓ��ڐ���e���{�S"�-}���v�؉W�6\�uO�����������m�MM�s�Ţ��!�G�+��*4��t2���߱�ڵ��J��xy3�7��h�V��!�zI}��[���˙�ˇN���X���_���$�Y� ��X��]JQ.�Wkn�M�7 ���#A:�2�ۑ��cdP�����y%���gg}�5�Y�締�~�O��ˁ*���gMO��t: BW�^%��i�,'h�-�*Åw���lؐn�T���ծ4�#�f�{Q���N�H[l�5��mt��QQ�8&��W-5A�����|��	ps5�F	V3��_�����Ŋ�#sҏ��.7��dx_�O�k|EmY?��D�eA���'8�s��VN��~ �#(����7��U����uFF�c����0���Pd���i8����rN���:=}���6�|�w�D�����g}XL8.�k�mj`	|�����$����o�l�+p�8��Ƶ�Y��A*�wl�\�����W��h���]�$D�/m��7o��J��+�����~״BH�����b������ݰ6�ê���J�i�H]PP���q�Y��38�8��h,k�L��]Rni���q;Wߵ8�V	$A�t�`��%g�X!
k�;R@O�Ii2�����(67rx�`�ONN��t͵�A
Fg=l�$)�":��輵��01�s�bq0�Z��%렺�����ZنC2&-4����m��/bŅdrhc|�1�q��}���"�ͧ��۴W�hԠu�.��j���?؅H�*�/@���ʇ<a����0%�(�ơ�$�x���y�6t=���Up?`��L�0!����`|{qO�'E�c�� �@��ذ�����U�Ki�M����l|�0�a�P���:)��i6m���24�a 6s��RO.���]�ge��G%Iz.�D5>CIViB�2�x��׮Iϣqpv�MII^A��lt���BT� ����-!0�uOeVJ0/�G(���#l���j)�Y��'�(F�|��:5�s X�}����L��3D�*�6�K�$�S`ƺ�o�HP�Z�Rx8����]s�����+M�*��96괎m�_�F@Q]�b�����+=^XF�ח剴��ؽ�Z�8��'��+/�����<�"��;�J�]�Ҫ|��bˁ��(��)Y8���\�_�Qml����_9�I���Q�� ��!��[���
�,]��4���I�II�H!d;t��s>B�Dx �\��y�85?�'�����S��}���E$��92����Q�_]��ٙ0��2 �DXP$ir���^�9�[d������r� �9�?T�]J�g��;|����ָ(:P����>s��B�l�ae؝�Jƥ�E��8S -2W:��4/��䕶l��VX�3���E'E�tfP�YP ���9y��i��{|�2��{@3"O5Hh�H��s� Pa���?CEGv|:�IIj0��n��A5Ho[�FpN�٩z7��S�����u�n+�ȞuW�ᦕ�Qi�)EVd�5��u����^[�ᦓ�-��bS"�&wJ���Ⲕ-=!!
j�ꉘ��
(�����g��01K�
K{8�Bwȓq11��>vʷ�%dh�EC%ʀ�]�?�L�s慇������ IY]#��|w�\��5��>?�	��Q���?��*G_I)~G����ޟ."��qm���4�q�y��F��-��Kԡ�9��z���E�m�g�k{9)es�X+�x`��@u8�]Q\!�7`gq�����b���+��3�kbpX�]�j����tK8~���U������9m�W,���?Ӧ���]��͙{�AA �}=[�][Ǉ�)K��+��kb��oƀ��6� �ÕX������`��I���܉Wv�� t�9W��9PҘ��`��ڂ���+C����b^�WŰ�`��"*"�c�}ϔr�U�|p��k_�ʔ���KJ�
a2gVq:D_n�lRg^�}= ��0�	9=����T�~vxj�i7|��8���O�8I�!a�<��e�t���	��[k�@�+6Ó����ɕ�R�) ���@�5��+*���Ϋ��O�hh~u��ǽ��߹�a�Ml����������k����$�����4�J��/��W�a'<f�5(�������U��
����o<�@����p����5 �塓�N��������m�9::&�Z000�bc���1qݎMEt��@�}N#�q�Dm��
z�Cz}n�`��;�N�~xx`�������x�O�ty=o��h-S̂tt��͍��������a-��͵!6#q���1��PPJ�yr�u�z�=��'*�=�F���=���/ �@B�|P1����u��r�Ɠ��k����ލ�m��X�X�swgCD��W �l[��,�$���;��0Yh�	�P�� �+�ν�P��AfYdD�z[R���w����Dĥ����D8s�����H���}u{���tF��ӿ�q��?��XYc�����ƣ�AԵ�~/A*B��ڨ��~H��ۙ�����Vv��	-1�1��y�;v�W؇�_6ަ���[�렍�m�Yq���c��|`]h-:�F�Y\�ӳ�z.���oOlޤ�!j�.\4m��_��]<�$�/���w���К�EY\��ݿ��`K�Wb���J�����5_��>�[�y�S%?4tN��O�'�rl��wȁ�I��z��t��>�
���m�CMA���D�D�0�������[�֝�U��=}\o?^m~�G-=�α���VN��zg`5 %%�gfg���[�;{u�nRu9-oĪ�Æ���`/<�a�~��?�"�u��x��x�B�i�Bw8����L�����"ؚ|�Z��X��o1�$���cy�G��B�)&Y���-"X�c ���:����G_�����v���u��7��j~0-�I�(��͙�i+��x�}l4d�� t�
~m�_/�UoZr��n�)*��gG��WH��?8@1p`�&q�Z���8#���\��&AO��nX%w:xL�� XH�.���V���!i��_���YSپpL5��������џH�T,���b���W������n�����B�|�|l�X�'�ru��#W �"-;<�+ƀ*ޘ����x*P��V���,��trw� P2�h�����+p�__�sd�4x P��V��q�֣�L��R^�Ύ}x���`o�P��e�%Ny5"������<�pm;�1dT|�8�E�ߝY���C�*o�7�+^�(�b�7[j��=98rbȘ[ �lh���k��]Mi�%7�j�D���*�Ҹ�x&���h`@%^��}S�:����ٟ�����B�9lz�	TE*Y0.{:{�6A�ؔOB�6�(�k�8���BY����UL��9�N���W����s���������!!!.7ä����`M!7��F��^�7ؓn�:e$x�P����o<��WB����&��(������w�un �����ȩў�A w���K�����~�g�(���z WTRRPVv*xsV��0�V�H�?�s/�@/ׯ�F�W弊�0�s��!Gs����t�(����,��C�2�̨T�oy%u8�gs-��!��c��T�0�}~)�u{��H���**�ͷ\>�ە������`�M�^�]\;���*RH��J�p��W�@�"��޵V D<)L:�ј�b�5 �KiHO[
���Џͽ~�&_�D4����}k��i�K�`�1��C��[s�JDj�<ؠ�]��'�΍�֠c�;���P�	�=C¤��)3����%z���HGL���n�C�T���L��@��dzlM~�������TP��E&_|���n���dv�)�� �d$���ڱ.jr�_ ��*�C��Q�W$��w����#OגKي�q� y�����r�Ke���q�)��V`�X�a��R)G�J6�1�C�	`ߣ��4h0��}��2y�3a8����P<h�·���Ʉ�i[��I�m�5$ឬ�$�hQ��GH�����P��mIۣ��cC޼�wm��	��
��x(���Y���X�\b���c�rֈ�D�'y?񾒷H�"ab��,]]�457�����F�Ǐ(���_i`�keRW����J;�ʰ��������p:{H��wn��a����~4( ��}��$�ibf5��z�{�$�Ȑ�X�:#_�������X��}�
�����퐷w��`�ZA�F#x�P�єaw��짓F��SZ3#	�z��9m�$��ѿ�*���S�f�T��6w��H�jѡdF�����B�y�ܞ�{8iA�g��L\�ţv�����D��A������f�n�q�����g��j�3ħ�Q�1w�c�� �����7d�x"($�I�E�����Vce��`��k�`��_w1|?� 0���ČH�ĸT��y`&[�h��OS\/;�	ck=w����4AB�\<S=cLa�Z�;wiMG>�2���Qe��Jٹ�+�Q�R�L/So�!����L�.y�����7�������{q	���R�\�6�h%*���z�h[G����B�Ky�e�2��~�ks���4{�����ʬ[$P��Њ$M} $g&�p�^�-��K��!��s�os��!��ʗ�dgu4���9��p�Ŵ�z��Y	['����t7\\�\k<�텓�/F���]�`���(An}#����tW�f:�B�ū/���v������G>g��q�����kL�qq7|ƌ�&<>]7B�5eL�xY���
^����XR30��%sߏ����0�8��f�tR�A�dNV�ۧ��JhKy��z>og��R-��N�C���7��uͽ4�����y30�� ���-omVq�_��v0qi�6�v�r2?�GÇ��Ie2$�!ɔ���UO(���ܻ�e��w�99dp�W��SL�
�����]0m�ug^�'�T*H�_��Q�@���r�ㄵ�, |�C�)`\p]e����ZQ�A����]���_ĊJJ_�����	�����)�~(���iw.+���u%N?q=��G��D�ŷ��iieVO���l��,^�P��4ٶ��R��h�,]��G��������k���ܲ����^-4�hЮ���-m')��*�������)2�.�u�W
�`�^f˙#J�S҄���*Ϛ��*9_��w����2xI`c����ӗZv�4kf���`���hRi�촦g
��ԨlY��=����Uk�Z�	W�ҫ���8�	@�rs֮\~��ٳ�"�,�z���7ؤ�(=�r�%����N��]����ً�rs�:O\,~����v%�ɞ Ĺ���vk�'��?���r�k~�Q0{�o��㿕[(��ݱ��ǖ^�S���hW,�X�=�H�L�{w��*�Mv{ZK�r 4�:���\����}�t�gyAG��کL��X�Q:.+	S���Zy{���D��i�i=��`�e
,�� G��{VEE�m�Hv�Xq��`$l��H։�����I�����Y�����ŀI'��٣�E�:�Ӏ�����4a�����\�'�q�,z��aZ+&8T	�=E��(0͒	����ҝ��j�A"t��t��	>���i_2f�Px,���sQ��\A�5�B��U��/Q�{��L�l�ܾq�#��YMs"K�Z9XԨ�(R� Wܺi�x���Ԕ�f#��@����%���/'��v~MW*�gP�7[�du� �B#p�tUkq�����ӓ�E�-�u� �<�I����"wꄚ���wH�o�������-H�=���6���˭�~��KX�YC�Әs�-���L�����������ґ�ys����ќ�zi��� �6j��P�*��Z�^��o#�K�}j<��;�x>,
=!��\M���FA�[�Z��ʔ�ǿ]��a�[����� t6ˁ�9��c�����[����Zk4�� �诋߈((`��eco�WG�����G|%��Uf�?�3�Le�)�` N�j�H̲�[���;=�����H�L�P�5�x��H	��3G�u	I	�c���IǢ/���Tm��	��ci$X��YK眜�v�EXʫS_�K���~�iv��LY�>u����3������s]��|���|�51�]8�b31��m��޲-�=�U��<�!c
5�O$��7ۣ�1��G��:�� 4\Q�w�' 7�"��ml���n]�;3_�B��[�4��M��6�sи�ɩ�OYz�'2Kx��Ơum˦���D���W��a�&n&����I�"-�3>]ͯ1l�ZQ[T��;3s���@�ǲ_��ٞOЖ2�X瘌�x�v�텢�,6���Cl&�3]S�{KQ��o�B��\������1�O�B�̘��i�úF�r�[S㐄z��q�*jj�)gbr�r��}@2����-wrҐZ�c�ȶr�;zE�}`>�52�������&��ЊX1@�㣢���_�V,b�SΨP�_��_���S�FfG+l9sUJ~s*�n�dD5�_ӛ�q���)� �x1=3������)G:��i�s`9�2�\��a�TD0��L��13�B_�ݔ�����n#!ێ�~a>�������U����<�,�ب_��Ul1T�-e��LjC̍����ioK�߶��b�H%���3���*yi PR4�����`tP�H����Y�nz☙�����@ǰ�x3L�N�����bͿXY�QNKiF�M��3:9꘮2Dݩ�f|#=3k/+?؏.��,[a5wz��Q�'s�
�j\��A�����]JUR;q�ą�6�����\��v6O��v�Ygى:==u�P&���A�hg�CS�}u�&%3%!McG�Y0G�p�Q=�S���<)� *���-3��~�d����#���S@\�i~J�v�pہ�Œ<9B����d0�k��H>�����%E���MSM�4���z[��|�#�(�����[Z�F�"�Lfp�|<���T��Ύ���_y&,W�pqÊ�����t.7�M�XZ�p��$���}�t�$�����0?�u�f��~��F������]W�g��a��mFoO�QW��"o��n߾}�_�U^o���U�ׇ�O���9�u�7	b6�q�S�O/̴����*�Oߜ�w/L+����ڀ�j��?���)��U�)�ů/Z/���q�����Xg999���/U���z���Ӳv������?ޑ�C�K�C9� Q4���5x/-7o�8����&�?Mm5�4�9��)��z���$��hG��lC����Uuue7�}���o}sљ��D��	���BN��Tⅳ����b0s��T$��d}����.P��gB�Ff�
�$�
H�?bXhnp	i��D��?�r�</z=vਫw�eKu��c4 �z22�V2�#�#Q���n��^C� ��s�|��m��,z���˞&��Z�Z~��� ��-O���q����8���h���{´?B�~4Y�o�w�m��8/�?�����{\S��,����݈�W]T�S�{�8�:�$%������=��B�Xr&O�"�;�S+Y�K���;��	�6�xw�rq0�)�V��w'���e!�6sV���|����P=����13�98Rґd�a�!����/n.z&��>��
q��`c__�U��*��ڠb;R}�����5z֛�֫�e�q	}Ǫ���J;�<��i-=�ʾ��m�{^��v&�{qk�TQ�[�,�x�	���Q�)paC4G�٦nMy�1��]ć������􀻞���]�P��f�p=]��>��R�Z]�x>?�N��u�N��sc��4�\�P���dq!ۼ��o���?�
�'��5���Y�*V�K{,��-f��A,��;���V�=�FIQn�B_/g3�z&������s3\��Q�6�A���r����+���U��Ҡ+!�������!^�
�?
����_E�P�vbO�v���V�p�g�$�lRXɺ����T�C@�����Р��M�A{�V�a-A�K�o�v�^J��&��l'f �$CF�zN�a��t7���p�3��G�׏'.����T&���{+<VR���Ʉ���J�]WB�cp��+W���B�E��칽�G����᧝ÓZ ��Y��p�Y��C2�p��/�r�D_�ي!I�����ǈ^�v�z^y�� E �r~I"�(�d�O�:��!��a.L5wpD�d�z��m�N�?aC���;�+�gex�7�ݳ�;����]9`��j~ˎ�c����СO�6h�J�M��:,:��S��ζ�~�w|a�mDā�z���J���¯������7��������惥���	�������kh����a���%d�^���tm\���Ҁ@���E�:�9���ßԩ$�-i)q ��������JĒ�tfJ�.=�r�XX-x��\>���~���C�uf��p��Wd@�5-��ԅ�"�|������ �{����ݽQ�q�z_2�t��5��`�n�O����rQ�@�ƹ�����'�þ�2��HTF�6e��M@��㳰E�(|�9p^ԯ�8e9�&cY��ѤK��$��,�eH�)�;��D>��BK+L�u����xq��G�e�Ȋ�Be��	��4�*�hf���x7��e�7��>Z��'@�_�Zj"���%bI��g'D��;kѪ��;�8�hV��	,�k�oo�j͐�3�w�a���@H�p��j�4�i�w�F��n��n�X��0�M��#��ŴNMQ��yq���H~�����P��|��b�頔�*�x;{�b�
��ln_�w͸z��	Ά�#Q�`]&w>'�����c�Ϲrg4Ȑ�|����U��yz�
�R4F�ё�j�t�����'ND`��:_s��b�+ED��ҫ�[�����h��ئL�텭6�.E�l��-{OG�C-g
�+��!_*D����G�W�7�������/Z�6���?��k������x�Y��g���L\L�Z%2D���*�������~!��]�˪/�fb���9��	��#�	~:�ӣL�\�?]jiii��O�͚#|f��N ܃��k�R	-">��N\r�Ѱ���z�ԛ�K�r0����рH�A���fّ��u�P��|�\�,�8��P�^��r�?�3٥ޫ�~���B%��p�>�;l���hJN�7~x|o{�7���-P̨	\	hhO���-R�HA��H<D��y����N��z+<�g��m��=���Y^����k�a%
�
\�ܕG'�}m���pA�_���22�9W��|%���L���=Z�˲��=�!����;<�Ma'���b�⟨����D�k�)!2����+�,�}L|� �ԙ�� ���|�����?�c����%�uCz�ܟ.���vOLH�mv�7Xt���Zl0����:�̌ʗH�;�+���e������4ȫ7�@����aH���l�ʘ;|��Ȟsv���+�Ŷ(`��:`WhO�!~�sss����c���J=�Q"�}:Cs�r�V¨�--��E�0)u�S��5�oj�+c�]~G�D�ѹ�#�T�y
\����c���v̱�uH��N{cb�|�;�۞���q�x��<)&K�p\���}�J�>lE���tNƆ�;LJ.��+%b�0Zس��q��� �F��󔯒m3U��}t�X���z��hZ{�V�����}���29!GOT��+"Q��С��#�]:�k�Z>�A�.}�@Ʋ���u�����;��S�s���V��s�<�i%�1�M���I�%⎑\��y-Z�O��*8ئ�*}�1�E��}QG�'V�VT�&�\�>Z|���W�n�RS�Y�:�M������4AAq}���Ɉ7�REo.��6��m�<+.N�Z��ĕ*Վ�zl��4U��]�A��P��7���v��\���o�%��?���֖��Me.�Y�?{�������f�#T�	��`_s�+;�s��(��1&i ����a�/'��j�>���أ�V,�g���C��Lds��L���[�:Iyr8��N���ZY�ʝ0H��.�ryޯC?>*�@���@�N�Hۛܽg�*����*�;�C��Z�9�7�7����?N�!_�d�ށ��}'�ԕgmS&5�]֋���ׇs�6z��cR*����E�V'ꯃ5EEşLsE4n���YH]�Xjq��W[
ƀ
@��P��7�Ϲ���@!`��.L�>Ԅ�G@Ų�NM�����,�c8��~q���a~~~0E�U^򻛛�8r�*�n�dFhI�{V�(m�gb��-��Ɲ��6.b���#$k��=�r|%w�������9�bzE(�On�t�hxd���M����"P���2\�m���sy
r��:���^/Ng��a9A0W����t_:��m�+�C	HȺ �+�q$1GN��)�,���}3\n����7#5j̿�zpO.�-)�1��"����q�A{��k�4�<nA���y��h�uU�ʨ�TBO��M�
�<龧�ǽ�^�h?�9�;�V�����
س�z��̘�K���}��[�eˈ�J�N�&�d���*�7T#B�7��l�|�X����@����W�W4���Ŝ#݁H��tF|
��Y��8u���Z�P����'��׳a����H���륜���़7��A� ��Gk�x�Qki]��U<|�/�oNCF*����;�@8��f�0����j�}���$6[���o��S33z�GVVVI��_��&y^�	���Ι��L��x�p���aP�$P���dum����QW��4���Ҷ)68)��lw2u��A��?@01۷���_ƘKae�#'$"��*6��,I�hJ���@xQ���z�V��w��=��Ð��e5\z�dK��k��ʴ���l��۶����ƙS���"�:�G�'ӧ� �\��<��� 
�r�:Xmd����������̖�E�Uei��?�z�&�����0�������ՇY�����R����X�}�5������,ߩ�ӱP	��T��:��+��	������;�~�mOU��y��5�g=*!�-��4z�c#�� )�Y
$�E*'�Re���al^+^��3K�5VbԿ�7�1mn�	�3��CBB�2������R��%پXo}zX���a������Ԙt���]ӞI�P`��A���.�ԛ�o��R?=co�ւX���-}hh�,XRB����[_�niiibn�'��}��E�C�������AXV���C�ǏXZRqq�ݼ��Ԫ􅀾:��Ć��TB6����qa6oX�?e]w8\[���Z��Ef"�%����È6z7��=� Q'��+J�̈��w��Ѣ�5����y����g���o�������mpz%iXޤhT C��1Eb>|-�)��yuǷ$�$���aٶ�;oL?f<�89�s�K~c��$=��8���ٵ�<{1L�R��|�bq����s �a;܀b�3��Vf�o�/��{,�O S���ᣉ��+�"��}70���8�sg?ȞD��`٠��������`mA��k�s�)cmk��ޅ���C�!�U6�}Cc�����5�5f��n�p�W�<Qk�(L���Ğ�拾�2��'���T���/�k�c����++����0ݲJ���N�0�����u�]�tA�����zF�}�����l�����a1��6
�"i;t�+[ �s�/kiiYz��v��JK'�$hJ{E��Hڀ[��3� Y�寽˾$�d?�Q���&���?�Ən�y�G9�W�{�Ah�p��3L�r���U���L�����[��@�G�jGw�<�@��Iº�V�[ fx(��6��+Sw����	��:��t�R��f�ӝ���s�b�C��!}�)׶�N���K���s�'�r�t�vk~ݍ��D�[��:ԣ���lj浾\�ND������[K�WZq�v�����$>g��}�<��(9�n��+��m|\�i�:�2�t�U�d�B��V��xe�J� Za�h��2��#�*��_��4-���B�5]���1�RٙE�0n�^�V.��o���Ŋ^]�B�ao�7��d�'I�����MW��	���19f9�]�H�^c�$ד�����Rj|c�����o?m�7z	����و��
������@9�h,{'=`�"L��Z�/U�z��u�G[۱ܻ��n��%m�yy�p��?������~��e�5!�MW��A"������޾dJ�z$m�cY�?Crbgk��݌�ŉ���k���	??+�X_�� �)�r��?�c��������&-jW�	CzBKB��"�a����@���`�;/��vr^q ��= "]��f�W"���DME��ѯ����7�o����u������$A[�4$��[K�%�K���d�䞈�V�2^�	&�Ϋz�����aO�3h��r��ٝ2��:dC^sx��6�ā�D�Y��4�A"M%�:�N��^40ֲ��#[�ܿ�+����Y�69t6w�X�V`=�ᰠ�UN��'g�u�;E�	_�E��~�@����?�����������>B�����8Lh�G&;mp�G�OM՛����V;�KrЏ�)s_7�}{���ￕB�7����P��1D�?���Wf�gr+Ɵ���~��(H��'����i��a\j���H���Oލr�Ƒ� WI�&(J�a׆�J�����mhʂ���+���T��I��&ݛ9�^G[|ڸ�����a�y�+�w�x��2m��	_��=FA�o�x�̓g��=g`-�Plr�?.��/_TC�U����kֹ>�c �37������*��V�y��v��Ïj�F���w_�8��)防O�GM������V��m�O{�Q��w�����B�,'�Re�A`:'�O���r�{��`,���w{�ϑ���(���;�M�"oi���FV�Q�$�/��3.�	p�1}Z�Z�lM�vX���è�^]Z}�tx�:�vr��R�~�Ǆm������|8~YYY಑tg�3���`�u��%k�f�s�~���ԬC�31i;9I��g?'���b��tM�5����C�����!4zER�_���T*������Mɼ���J__��{S?�6��D�Ӌh�k�*3��μ������#Y��Q��0����lD��iSl�#�o�:K^mzY��|����7+P�PK� ���������wi(���l�?ddU��R=7��cڈ/1r��+]V*��>Ƌs�7*���:H�-�S����KmgꍣΊe7���G2�J�
_��'��ѕ3�wߓۀ����HK}��իӾ�VA4u��B$��e�ϔ�K��>Vy@cA>K
��R��ۡ�{�I�T^p��d�րb�w�&�TA�\O\�BMy��LPF'�l��$]���S��f�Ew�$*
6+F�j;��Z�e6�����I�_i9�)��v#�*� exf�d����b���������ʎ��^B3T���[�v�y���Q�B��K��q>+}�W7�����?���+D{�7���u���[,���"4�.���#��H
��s1;3�m��IyI0X��h��E]7,lru��h`�L/L��p���p��7�4��؏��̊ղ�ߓK�e�,o`ԭ�eA��@�%&QE�9<�Ӳ����ص�ai��P�e_s�G�O�BG��n��X�ӄ�:���[�bX1.LK灓j5�qgVf�Jw��x���;
���?L#_e]@|��oـ5wc��j����%�+�N8Q�����:wR��v��S���	���TT{$:Sة̆����u~�}��8��u�w,��v���şw4��^i  �/��(j	��"H3����o^�>��t�������+�J�j���̹�XY�sXJi[�����o&�!�D��L~*3�c�.Yn�s���E�.�����}�LT���;�@_���wTz�����
�q��YO��7�9���#b([Ξ�9"6Y��8�/!���l�<�l�!M;M3v�	�����3�_����9ܾ�` ��ϻ��6�%��/X�9@�����^��LhjR�A"E%%i����M@?.v[LJf��54VT0III������S ��>�DOnn��2�-���W#�ĢMdV{|Hc��x����-`hQ�e���I��P�vz��e�%xlf<˘Y1��Nm]����^�ݚ*��)rs���h�Z���LL
���q2�@��vZ�g�"S4��:θ"-��0�'PdMbp΂�r6����	�Y,�meN���I�+SE�?a��ٮ���9	|$�y�yߪ��WB\�h̄ʫ=�9x-��X�F1��Ԋ��Z�vk��/��}�2Nh´�pv,��;�IV��<8_uX��r��_�Nl���:�^lb�������4��C������
���޳YT���B���a�[��Ү6P�˹��xs挠�r�i�vP^�}%�M0�fg��g_��+Rr�>CԤN�,�-�^�F��@���t�����ڔzC[F�Ȋf-/t���GQ��<����"�Y���j���m����ꨭ���^85VE<5>P3<L�y��4��o�ْ̧�M�4�������$��[ں�=����D]}�MG�m���'O�Η�ѫ)��� y�7��/z5tth��^�l<���D�՗�3*W�������8��`�6@��P!��"�ޙ���z�`H��H]ݚB;#(�{��,�n�h^�E�\�ʠ8�U|�Qc��%�*�����d�kZB�#|� ��<`��!x�
ryg$R�S�'�
á�I"��`](es��ς	�I��u7H���X�
�"t�*�`mi�����̯Y�δ��UH8TMM->))6%����zn~~bj*fr�ɗ�;�ǒ� �+'`@+4Ti(N�v��/o��[l9�����]zt}�:� ;X��j�/�–+�-Xn��T*� "b�e�ub>=L�U�jTK���C�&ߧX��q�&�IE+mŅ���m7:Vg2~��	��)��� )M�L�ᖀ�+����y3��0�����z�7���V�ma���/�5���7bz����y)b)�H��H�+08P�"]�~s!�;% ʀ|W��q�%E@s-�����?~s���ӟ4�=pc���O .�@޸р��L��T�h݈��1���3p����v�,f[�H:@�N+�s!��*�ס�x�d�
#�������T�Hy��
��e�y������RE �E��ʸ���o����o�E4��@�V]�Q�U��`����%���o�B/����r�ʠ)H�f��Z��6�Fd�`�1�t<�6���a�� PK   F�Xࢳh� � /   images/554ca8bb-9ffd-49bd-8b27-eeb836a64b12.png\�X���=�PRJw#�t���4R��Hw*-- �!��-�%�H��7���s����.��f�=k��֞!T��"�BZJ\AX�@ঐ��O�j�r�?�E�U����q�7���GG�����B����靆�[S'W���+��'+G#;f[��#"�"-�V�-�p�U�������\��q?"�e)j���wJK_Q���4mj4�$I{{4�
��5�gg>�-~����S��
y�CMƷh��!��,�#��f8j�cϣ�"!����0~=�g�W�O��'=t�ǌ'�g�j��H���mX�ߠ�Z&�D�O��[��[��Ʌ-Pvh��q���hGy)��>��%�|�����~վ�8d��Xt�x�bgZ,���T��e9>�����?�|̈́�"�zNX빟z��x��L=6-�.|;�H�0q��?��|�p���9��e�ϣ�Cv�~.��!�o����0IP����o_��|�N��N.�؜D4K�����vr?r��i�?O��B��B�a P��ۅ�g���g�!�n��Z�g����H�x�i	�֑�Z:�D����?H1`�[pR��D�˲��c�k��q�g�lwC�=��$��y���`��sDVT߱c��7�% ������.�Ň�K��s���&"�Y�@��A<����7Nv��{��Lr�@��)/�?�UA&og����E�i�|˽�Ӂl@J�W;��*
� �1�[_J�i?\�[������r�3���gi*F)��yދ����BV�?�5�U���fv{V�#_o �@2`YM���8���" hpf�x��qv���a`5���:�TS�hG�"��$�3�>�_)$����Goo�����cdk���z���!����H��0���A'
q��D4?�pR�ٗo�7_�`�E�򋴃�(QD����!V�Ui���l��C����YM���vH"��p�����v���q�)?�%�dY��?��8�y��<��
��3�h���D��?��Ly�cEm�
ڠP�h��xVAԾc����07�>?O���VQ]���Ȩob�����������sךߐ�\ؗ����V2���ndc#?D�ޞMFVVIQ�ĕ��Q��Ghbb":6�kn����������>��h|����	����U�Vn�g�݃1���s$���b��	QPQ�F��VU�|���V/Y���
�6K�U�9�lF<<�ݹJ*~�](��y��Ӄ���<6;��I2==-%/�NS�:����9���ޗ,,
���?����F��><�bdd���Eb�;SViii5���XBn~�zO~HD�;//����x�`�zX}"�&L��Z��Db��6
e2����g����/�����D�b醆�w��='�hr=~���W��slkw��]�ܹ~[��ث_?���|�����j�R�/y^^�\p��;$�&pO$�L@���O?��?��:/o�?^����76��~[j����z������tѶ���9r/���e�Kr�;'$$truTW���Ĕ�&��&@���e�3B���^g�"!!�l�` ���3.�Ѐo^��8�2�3��pgee�����������SNnnXj�&�w;}�5,,	-��{@Կ�@䏈��G��\XX Ly"77�>����zE�C��,L.	"�g��"[<?�S"�8�����',,�X�:K�̃����e���Hڛ��
�M�r���],���V`�Q_��
����\p����F�T>�g���cgZH��E�}���N#��5vO$����AW���D67V^�I����nq�E���Ͳ�?�g$###x���I��g��4R������j����B�ݻ������8��x�q)��A�(@n�!g%�urr����K�0��k�ѯ���u�����qrb�- ��.��ӧ��L
xD��`4���EEE��� ��W1���m��ڟC� �<
��K?�0gĪԌ7:[�u�����h�M�n󍊥S0M	5�'�oְ�&0'rY��*�?�����'(�k�ps�$��������"�g �HB��h�$D����l6���Xۈ��4��j[�qq�+�z��l&..YT���D	VLLL.C�4++�|��krͼ����b��(Mk"$�7� �R��1�ǉB~|z���~��aK��͍��}Ulr�W�F+��nO�����nq���R6�#�_��X�'���x]�Y��i��,���F��� ��R~��U���+���\�94;�GF$�|�2F�����,�Pт���PQQ544�'&Ύ�OM�}���TR��L��%33�o��G<::���T`������g'�������\�sO���o�G�������L�[�qf���4�͑��W����[�����u[:km�6�1�ff�I�p��A溜(�	i���W����_�$�d��0������		����ݿ���MKI)�s���+���|e�ź���_�ø�� �N�]W��C���?�[��s��#ߗ/_���"h���*++���nԏh��pUUUQRfgf��n�J5;��P��ӡl>׼X�'���Ů���,Q7���E2�L=G������E�=��ˠ��p�l`@y���������������z���?�Yb�N�s���W���\!qqq����58ҁE�		����wVW���Սz�	��Ǖ���=��o6л{z(�� R2Qb8�)�g-~�,*Q�i�`����`��l��tRA������!�H��P0fA�D��nYI��@xY�.���ǳ'���ꆲſɗE��O�Bq��l*_���p������\Ԫxn׷oaf�t���
�p���܏�-\x��SʯA@J<;���%����vpW"�������.��鑕�Mi�<����L����/��F�K����pXUk�����e>���/�u�T�nw"/̯ǐ��wZ[G��tK��MIQG�4��VY����XV����T�R�D׿���dˈ'�j2���ťV�nkk��l2�:������)CQ���f���Rl�{��������?��]]��},��"����6��Ы���Mj^���N� KKKxP������$''G�$�ɜ���k�����(#ݚ����X�*C/9�����RJyy��@,�(..2�#("ZZ)�}��vv���Rvǿ�V�����>�s<�V����~È0D���%��8=g]��7����W����7� 0@���IIl����I��H U��j� ��UUi�V:W=P�����m�|0���z]v�(&&%�u���d�i_��0�m��<{x��>��_��ފ�@6�ԥ���1�t*�p�b����χ�����X���Li�h�(�3qqx4^��8��_Y҇��88�Uf@t��t��55<:��J��Gܨ��YS#�sp��lv!�GT�[��������\6:V=��H3_������/]�suu53�HQLL�ϠpeHQ:�c�i��{����%))It;$2��蘘��S;�v^Ey�@ t�	��P�Y�2����Zo�Q�j�/,�1�Qc ��Y�:��B�U�O���d����Ǉ���M��B߸ ��ʛ�p�cL}a������8������� ��tAA���;�A�"EM���uv����$��<.3���lf#$�I�q�H3�6(�C����כ���1!O�\�f,����"j.�֛U���=n��p�,�)�����Q���c��H���1�$����-I޸<�֗#�)�cT]�W�����I��/���B�<s6ړ��F]6��;�ӥ��t��FNc�ں���r�{BВ�w\2CE��_;����ߗu��#m�E�5���~�k��SV��5�@% @�Y�hchU��:��Z���k��	����SPl��U,��$u�������h�/���*�ZJH�mL`9>P5��w�*j+G����-n�B��%:^'���G[��ѱ�*��A���Ԕ
<���r�i¿�&�eX����µ������W���D>WDO�th�B�����S C"�>>x�1�����c��J������l�ke]�$_	���5�Js ��� ^�K�r���/�KD7��F�����u5h@u�M���iry1�//���]�/~��<	M�R���$�5qO���t����<����Ah��O �"P!x���s��=x��6�Veqݍ�7^0?�F�&G�λ�~���Tn1���p?ߦ��T)�{$��r��\�;���&���4H��Ɔ@`N�c2�1�gH��Ի�xI����|!N��� =�6��)߾})ժ{��%l||�1C`�̷,���+�+�z~46z4{'Dm�YS�0���"�ᐖ���J�֚�V>-��������$|w׼!�b
�ĐI^�G�V�������91 )���HME����瓸n��c=1�ng���[��3-��d�Am�f�R��!����cE��mf|ǝ��>(>|hG���	��J��������^|�ʩQ��F���[W�:vP�p>�yc�ꚰ�x�����
�����~9TG�j۝�+��擃dOߥ��QQ�1��N������oV%�k]�V�Nȱ��&�qA��+)G��2�ㄑ�u���Ə%��������IsQ����&����˃�:�M]C��e#L�yy�m߼Z!{`ߺ6���Xb�倠���Ǭ�q����4��(\�V���v'�&�	���F�c�c����s��J�-��~ Y��;�VPyۣ槁��F��a^���_�.x�v����Ӗ�~w�r��������r���)�U�6�p��,(�=�lF�jΔBBd�?v�܏���$��sf]���i��y�)���+.C���DżuC8!)i�ؘbn^� gdC!&���X����má�LZ����sP�7q΍e[���о�~������j�}g�7�-�#���s|:b�$�z�?�#Og����S����zݰ9G�p
5HxxA�<�%%r�����9�;j����1E��R�C���,&[���@+��\^��z���$
y�򁱌U2Y���z_%,���W+��n"�}��]���U�yC��0<�δ7��d�]�9F��^�BkK�����XmW�֮=��Nnh,��V�T��'���n�*��P'��ǳ`�ײ�u�u|��v����K�"������4�\��'��
d��/.�O��<ߠ6t��tw�ׁ7��7�mGUT��y3D2�Fx����df�i�9���`�ɺ����b�X���3�hR���h��֐=P��o�����</g�$�<��r_3X����.�G.��Wj$����
�c��'� #�"I:7�����F��ơy�;G��v�q.�����`f�	����CB���Z;���o��A嬴�D���M�A~φ/]1
yp�q�'d�Gt�#�ׂ���������>޷9l���%��u���#�{��)���%��DA�ّ�*N��e�\P���
�=�g*os�t:�Ф:���U��v����N[�HE]G^^����4  ��f��Ya�a�'�co��K��+�(����T��z}��Ra�&j�Ҫ������y���T� �&���c����#���sq�!�qr���l�UT�����Q$� �`��}����Yb�����G��XA� ����r��mk� H�ݽ�گ����]�ߎ��a�Z�X��g�&ᡠ�6s�g�Xt�	�ǿ(����AA��*�#�TRR�����F-,h��uK���s����6+E��D����<�Ź7s\y�����&f��p�{�����ūW����$WQ�-o:��.}�U����iy�ye��umV�����܇I�bVf&��2���~�;i N@���Ɛ1�j������Dw�kw��Q�� lֵ�l>���u�Y�$C���4�p�r��>���F 0�¾�����|�fJ>���c�����a�ʙ;�H (����&�w�P�������=�n<�"2!�'�ѱ1���NֺL�@%bP/�.�i�~�6�Z[na�v��̒��~��ES����Ng�'))I�� 
l����A�T^̝ь�S��"[h�������?��YuEs���t4�i�700ꭊJ\����a��Qu��o���<DPVb돣)�N U��J�fL��H��>���m�`Pz���������]������L��-��GG~o�EV�Ə�T坝�fl�>�T�S���ޮ��eot>������XXX��}�VY�
��/�b���~[N���x���v��4�u9�4`�J����])R���. J+|�|
���!:0��H�@�������2e�[swvu�9�$�6 ���>�+�:�w�)�r",n��C��1KC����Έ�IX�U?�����?<�$?���A�vE�y��A���7������9�s?���B����ִ��HO�*vVqΰ=��[L��>��c�Ɋ�˳��"��(��8Y}�SX�P��F"xjIL(�h��+?9�m�g�=4��C$�!��X�`�t��b���}H,��1��i�"ԏ�*�`w�@�_��@.z=��@�r2�=m�6���O�lT�k�_y�R���8�ʎ����� �Ry�a��]ik�Ji���|����̝E^Sr2���Hꫫ��������G�n-���J+X�b71��OwJ�VGCC�w>��#�)(@�7��:���L���i8֒`ۑ�B >H���p+O8��ҳ���ggo�8��t��������VŨ���H�L��$ �Z�g9����?�l��(G)ih�������l�}�k��Vm�����8�o�����篃D�C�𛎡�pߧk_vc����&���eR(�y^1�z�q�݇N��T���xs3 ,�5��SYJ�#j�yX�����/����Q�����0���a����$2��٦��p�G|P�4�}�j7U�:�5�j�_�u﫫�s��P�yC|������?�bbb�m>:E�c��o�o-��ט� ��p[nN���k� �r�l�B�_�/��3��d��-��g-XA_����A�u}�4�tJ˄����.���� ""n�88|)/gy��O3���IF�{�ij��͂��� 3&%�د����&��20"�դA�UnԯQ㝉���@Hl\��WUUM�KH������Q+��`]$Ok���{���#��T�_���Kc�U����c�����:ۡ���>D ��=.�T��!~�f��g1dׁD����6���҈�
F�cY�Q��S����  �O?�V��±�J�"$ѓ�b?^�x�%�F1"�P.$�8�����NN�u�����,9ϸm�V�Yn���>�5���-������pgۦ�K���N��GF���~��9���u`�k�>����Od���C:|QӪr��cTIt��7^���\&:E�Z[���zw(���tk�����Eb)n����`�C0}�S�%܃م]�����s:���	L�6�^��G8q�x�<���j?��?�b��m�H��R�b�ٙSJ�Kk����2� :P�b����^��9����Y��
H�ݑ��W��W
�B>�f�uhW0��.�k\w�O�ڑi�����e���^�������I 02��)�ʗ�ee��hd�.�@�3&��%�Ѵ�~��-�����X�����5�Ĝ[R�/�T���� (E���@��#�H����И%Wt��Qz(���</��Cf�h���!��x#=3?���<ؿ%O��4)������8*�b�!tr!qee,��kR��`�'''��^�}!!%��T�~���V!2!/ ��|�$�߉���ܕ��ƞ,�2��-OΜi	�`cck�x�B� E��A/���X[��{vy�����HG�oNk�?�[l��u^�|�H�cKK$���Z�<>��dE.���-\��Ϛ�V�.�?���eS��a�L"�ת+_����ï�u����it�D^4]���*��@6,�ܰxx)���kV�M���}�����LL�C,mR��J�)��j�ye����	EC��Y99�ml�&�̟3'�
e(�/ S���<�|��cݔQW'n[�y@���^����h9o������h�����0���J8H�:������Ң���=�QxXf��pP��������=6
;^���L:?;��"��Z��_�`:'55<"It���;_:y�VݧP�֤BL�T��S�TQ�0��"k��=���Y�G����Дq��i2Ta��]x�u����Ku������,��6-'r�5�|Z�6())����,������NV%�.&4�L�}[�vw��l+SRR��c���_���NL(W^'`B�I ��	y�e�V����Pd� t^www ���wF�o�L�Z���Bo�&����@xl�KI�h�|�#B;�о��UPX�_�[�����DE���	�tj*I�NMUUW<����>�E*K�=(��4̠�����fKKK#!!ez� ���x�1 �(�+�᳈Mq��['5k��W�XZ�i�W���=QS�����4opU��ʍ��Y�d=�����B��TG))$���LLL�;Eee�~0p��Y�	�l5t;[,>C|Ԯr��v���>V�����ô�#���IĮDY����F�`��w�;uV�h��z	��_b �������*�����k�T�V3���~�fp` ;G�olLLJg.w ��..���m���F��;;:�98��ϛ#F�A�M��ޤd���R{D�i&�_�lB��h:�%=}{��ߓ��*��=U�u�jsL�ù���0|Û�5�$ɘ���<"b@����%��>��%��b�[x�Wq=�ѥ�;��|u;�5v�Y.]�a�HUUu�7([��qX���������X���4��Z{�< ��`k0^����� o���Q͂lN����4B=��z��E�i1��n�EI���W��ФWT`���ڦ��6Q����6Q(a�%dNF�;���{�zd%o=:<�.CȻ�}���~Tٝ�\㦠��Ɏ�UJ�f-��oߠ���2���{)H��X�4gF��_lk�� ��^|��������}{�HF��ۯZ6��r��5p��K����^����D���@Cջ��<ޚ�����[X�rYͬ�k�z5���p�d�ol���Ȑ��F����bӭ���ݫ��.֡�3kcx�m�dgW.���-�������v}��?��x�r����ɷ�Ը$$��?�d;9?�f�Y�`s�#�M����,0�P��,�Ŧ���c�9��ez�ۊ����g@�]�����O T�WGk�{|�}���Ng=����p9�f��zg�๹9�Q�J��2��	U��\�c��u��C�\Fr2T�Qp|8v����;Z�����~��������f)�e@p0�`��a7�Ĺ^��\�W�B�N�����©���	C=ߙ��f��)�/�++L�����G�}�&gfz��2@oA$�&�9���
<��2S �Vs��*����N�x������2��ˊ���U��6�NH�+m� ��TW��2}��_��<ӆ��aL� e���%s�����l_`�Yfn���	x>���w3�;W(++����H��� n�3Q(bRwIbJ�(
68�N�������c6�~��O��3�T���7���^)		
`�/���ɗ��JK�m�y�-�r�+����Z�N�����]�rY���E�"�l#/�n>]?��bie�)��q�rMa�i+;���z!!!@�o����@Z�2C�^����4*`��������s6������U�=.���c����rwo���~�X�f3V���2�=��Q�|�R���O�B���^ù
z�3mYT#�FsN�:�}��ٰ�ck�p�-5�T|f�� d�?a�mjɬ&5~	��p��C�o� �Y�ZTЦ[�НԺ0�'��} ����"�C��k]#���1�HQ�L�N�Rv�t]z-�o���:o=�:�O!��'Њ�����)Ѭ�Y;N«���8���C%�>X��;c7�ɲ�6�!u�E#����Y-�W�zws�a"C,wz�%�sO �~�D�,��5���N��n�h>wx�Eyپ��I3��|;T�Gs3���^ �
�=e�jd���"�ҡ�>��NP	����r��z���a� ����^���,1�������� x����!����ߋ&�mZi���j�a�o�V�K8D4����\5&2<��f����YԜC�L�����z~�5Z��K{�p��N1��V�Տy0� N�B�s��l�s�����Ӈ�����c���Њg���Txu�'&q����3����b�b��DGcX�RcM��w����wP��f��I��6����\�Ld�����b���ؐs0k�x���z|3p�_m�������\��ׅ���e}��_;<7�
Z�)�g���L�)����tAh3�OVVz=��!x����v%R�X� ����N�Ύ���, z�'I�
�yq ���J�p2A��SPH�ޓ�(�/cu�����p��PS�����<Vg�W���ա�wݝ�[sS�So���=oj>>945��*UΡG����ʗ�'����>��3@d�����ND�_�5	���s��UV�����xj�ZtQU<_t����K;zy}-	m�1LYZZ����"�&���ڟ.f�s��[��ͥ���npx���N��U>#T����4�O�>�TϬoh�����ko��E�VA�g��(D]uuD==��O��4���{{{��{4Y&UEEE��bRy�EK* +��ɥp�����LwO$��S�Q_�D�N�&�a	����x�����9�5���B>���,�����d奥�%(�B�ˋ�n`�u5�=8�g�7OS�Z<PX��xz�qR�� Sn�������S�g�g�/Ml &O�UIE��ֶ�������!�_��=�0�\��P�����i���E�6(�hҩ���}n(����QI����b��U$�4k�o�%���=�߇�uP�����i��#*�:�5>��Dp�E����))}T����!᣺z³V
1�Z~$�uɝ�t�7�Y��z��8��k���8Z�R`�[T��Dƶ�F�d���~��Rj	I�Ht�dt����UT[�����J�^"�z��G󭗷�;�p����(�g������v�@�---�l��P���)1�M'U�����ݜd}˹��E�����_�ڑ4l���d"���4ae�w䶞�Pv��s����(��E��ϟ���-��猇���Cϫ%"I^�� ##kT��A�:^��������@���al�3���뛭~sQ�U��=�K���I�555��.Q���<���5\o��t>10�2���*(,�TW��!�ׯb�p�^���Z�sH���jy�亷�٣�k���P�=F��O>kD�Ȫ���Ҭ��$�YE��	����`lQ3�p����r�Jؑ�ѕ��"U~'$�^�K�,t?�0���j~ ����XP` �x{�gmm-��jo�/"�E�!�����&��Q���=pѣ�GIE}6���F�� �N��#Z�gO��$!�-�40#�Ŷ�����ǋ7�����˓��Ri���)	(?vv�k���x�͛��������-|gjJ��H�Fe�g���ـ?~��}N�Ù�@}}��r���>�>�#�f�n��sgU�Q_�������A�F�2�Iqjb��	=Mcx
8\+����������-��|\��@Y|<.��>~�	6��ٙ��W�
[��6��^`{� ��f>FQ�R	>���!����鳲�Z���:NV��R�!1��`2a$6�n�`���^�����B���k�$a���9����f<��4�Y,.�<8GY1S�S}P��y��7�v�n�Bi�v�{�s��pO�Y���a�p&&99N&���eD���>l�t`g���#����VS�P��!�Y��/*�<PqI��6�M)�����W�͇4��L:v��p��t	�(�z����##s�����XW��tC�ի�o�s�?�!�����щ�^�Bѣ}���9��g�ղ-��P���"��d`�����l	��������X����V/B�'9|���C��|�pkڽ�----c33�O��h`�3���5�+-#[���w�5"��
g�����������tttY��(((�#��>f&� ����� F��A/�s��T��9� ~@}HŃ�ᇓ8��|#�~2�6k���~�p����f��&ZI0o���RP��Oo�#���A-��A�"�^Aڂ�M@h���d6�3[9_L�x	�T���{�㦰��f�%�W��o߿�����c�M� v�&�ף��0�F�E���`�����3�dnb�4��x!��z�*���=i�dY�6���j����������y$ȋ���&)y�x.m�B��G�"��Fq�H���
6Cww7�C4����������N������6B{a^��׾*�&֖��{:O���s�]���ru��~FzMcCkֆ��@�a��5S��e���(��4��Ж�˟iNiid~�Cz�ݗK����D��zm>�/_�$H�0�D���~���r�+�hk�v�5����';;;�DlY�����*Phdf�u�T]�{�f{1W���5�0���FL\��n����ͯ�Oy�K��z<>�}�9�"���x�~g�����~�`kk���杻{Ô:'R��IQa!�����Mu��E;P��l���H�GF���uQb(�+�&�^�e�N�/'�^�m�~��RDd��Yv���Y�9��Ϗ�8ѡ����-��~&�lbxQYᖉ1N���ԑ՟���/M���҉��p��f˪�^�UrW)V�Mb������4���{�ƿ�����u��/��P=x��!�"� ц���ٙ욤�q�Ս�5��::J9\I�fU5�f��5�;��,��R�:�z&�3���u�T�c�@N�y0��%|/k?07�!|�<-|�p�5,1R���1��wm����*�h+�--���j�&mhj2��i�KQ2�M��4�Hyq�9�K�;A����AJZzB�8Vi�'�d������I�]6�%��=�Y���6�7E����y�<��M>�x^s�9SQQ%���?�H��%0���n�mff�pi''&��]ej�'����p�~*�r{�NO�?&&�n`0"33�6��v���S��V�-�٤!����j�9,����9ׅ?I!��.�=e�?|O/ن�m��6K	�m�V�3������]j8O�eV|NNN^(�,3�%�Q����1R�O�-FVVŢ���ь(:�tN�ߛ���5��YlA}Ⱥ?�#|�����rL���G�/��XfҘ�W�h��L13���f�=j�f��&i_�|�;��q+򺻽5�{�..�F}h���_'j�Գjj�c޹�Տm�F���-:��BQ�2%���?�$.?T�OA�i	UX�h90��j!ss�bSRwg�N�GFGv��y]mC6��`�������Ҫ�����|{X>2'//أ��E��24lZ9{�s�����.S�Ţ�����a��Y񂓔��SQQџ*Pr{zl�?��p�6�i�~8��r]����q�M��ؘ�e^!�1�s>�r�_�i���G_u����ԟ��v���&u`F�xݰ=�rzc5[_��9�;D�ia�=;�n��]��o�㤗���}��K�]����pJ;XD�;v�[]�0���f��z4�	﯊�"��B���,��2���wu�!�����I��?yE�����Y|feuٌ*���+׿��hF�a|L㵇�4��������'��CI�#��ZCY�>̱C/��Դ�S�E����E[{`�A��ϑt�r���۝͛��0}{{�,8����"..����i�]��I�ٙ�V>���P�ܼ��R�^��>R�Z|��W�APP�_Α�����fN���5����R0����!-ϵiU���EGE݇����\{d[W��p�#AaC���Y�>j���ҍc����-���6���}���;����t�>hd��z�vY��C� �f�d&j��bb-sެXpa5���U�����}՛\\�N(��^�Y޲��L:�1�����6M�y�Tͯ�i��,c�>}�!e�Z�I�}��B*T�P��G_�ʄY��!�;1ip18�񎞉	���,W:����O$P��viqk}�B���g���1h/�͘b���*�������!�(���7��t ��ZCj���РO�S	-�&}��-�����DBFF�ENL��ʮ=^X ��]Sէ�j���3e:վNN�*)�X����j�_erWEq{hZM��'��;>�!���36��$}3��'�ERk@m�#���d����:��o���u���l��/�,x�v�(���ج�?�:�Q쳮#+�Z��"��t����z�jp��!���B���	C��`��b'�Ə�P��NY�tt�4h��K�+���+.�A���������u�,��t~Z��{�����)Mڼ��������Fw��"��/h��>?h�;��3`�PCK���*\�z�.+7�)�������HH~YY��V����ƌ�-��ԢL�nQC���&`�����Uז�P�8mߠ�U7+��z�Ņx��Z0��IdE�j�="b��qoUEE;�ʀǥ��`��|�e�d>�σ�t�I��N7q')��2��)((����兪�-�F��˩`����\j�Vv��DOH��S���O�Ϋe��Z/�|uQe��ͩC7�'ǲ������r����McF�F���:�������YI��G���!8�
w�v�$��ҩ�ZM.Ld�>�g$�:��҅�#l�r_�6�k���,;��	.Y�� 3y�j�<BE��Z�풿J~�8|����{��۹�Z�]���ʴ_��4��1lFkh���)�205�u��\��d*R,��z9ѓ���q �����Q ^�%��f#�1S�D5������M6���=��Sd��OZ���L����H�X�F���K�~q{�Y��$��.AtY^�Ցu��p�f�.����e��(]�@���4L�|��-t�����MD];�Vp5�Am]u]w�8� Vz��@GJ\I�{�*��q[������-�^��^K����"��b�ur'|u�J�s�w��T���b`i������"�����ʖ�/N���7:g;�.��[t���$�nhh��jC�{`����
���Y},��~wY5�B�}�B��f���zkߋҦQ�Hy�Em�'���{L��j����M�����FõNS��f#QQ��_�Ԅ���uS1�񕞁ð)+�dP���8u�3!���7�5V��L׊�[;����,�� ��E�������[#R^���&�9����ew�)�"g�݇�D�R	�M����7�濺�S<���虘�1w{�P��=�K{㺉GN)޲��G%��Ǻ��?l&�i���	���*�IZ���&�D�G">�����
\	�G7~�,�/�?�p��20`��̢Z��}��`��rvN,��>s��,����z����)�y$�xKӄ�R
\bVɀJ����sD�F[LRRR�BtDaaa��|U�Ʃx:O������KY7��ԓu����>� I9�ɼ��O&�I7P�rT������غ.�ZE(�K>V)�2��.Vg8�������	�� R�O������iA���RdFF��ާ�-c�)����k081 ����+m����!YM�#"m��ڭB���'�$�]���Ņ���ɉ��������|�"��ׇ��S��\�z޵� ����
Y�UXy�
T5����i�[0D�3v�@17����ʛ$��Vo6�M�лf�[,�w�0�Nȶ�6؝Ģ}M��E���T�ʧ��!jN#F<�7W��S��s3	�d<�
v;P�z9���>���eXO'���1�ӯ��ڢ~;�N"�K��z��:�R��� �]����g?Acdy��	jS�Թ6+�Ӷˍ��5]�_?:4Z��;��+K�$�nb�<u��/�n����ݬ��P%m5�3 ����q罹U�yzoo���=֐g�y�	D��kv��R�����;FG�Ǎ�ȅg��?ɪt.�� ())���#��>'&&�쭮�|knN����TX),�E�4-==�[f@�UzAF� �ѧ��_��/4��3m��C�?> ---5�ā�]I131�js�i� �����wr�^zT�=�ZXR�{A�h���������`��ߍ#m�x����z�?�Rcl���$�O���em�J{�KK+�#�^�J�MD1��-W�4~��,�K� �Ï
�2����g�eȮ�~&rP8#;E��];����W27��B�k=ۏ�v��,�����+��KQ�SϦ͸�������j�u�S�@�Z>"����Ïl��?*�J5i�U���i�/FA$3�]K��}Q �V��=;������_^�IN�� ��t^J Y��04��.��X\$u��q�� �w�$��"�����T:��Ď�MLL�?,�Z����f8�+]PXhq��2TW���&@�o@s�@C�8�8���=��%q���4u^����T>l��X��u�z�4��Z�FH�6N13.��E�j.�N����`Z�qZ^���ΦjO{v��Z�y����=W��|=>H�KV��`1Cij�k�2��=��k3�tѻ����RR!cZ�OgOsM�'E���+I��{-"X�~���Y��z���[�8J0TH!~*�_�`���H��Ś�b���k�"�g62��gf�Sh�\h�s�Γ�x��4�e�����rց�S�m��R����tbr���l�δ⊷k���1zm3q�M�Lw�R�t�����������1A�Nii	A�����n�n�H�;��������<��9��=ל�g�������5)��F��R	�Y��6y�@�O[o��``�l�Pn�(�.�*�w����v��*����5��a�+V�is��ժ.�����b�_�M��㿣?�,��爛�O� z�D	P21�'2�x�!�'��ܑ�^���n�/�'���0+<�y�O�n�y�;Sw��$�𮁹��!�m��(��n��k��ha҂jj��{a1<ϲTU���p��ez_�m�+�"�D��{̈́��*��ã�j�+����{,8����j_Ɔ��eN�Z�[��`��ͅ�?l����}�P�DD���~H���1_���"%��z*��x4
'���9������eV�����I
�-���$��0�ԋ���B7���V3��ӔF�}��v���h>�O����uy�ᕈ�����坝p���H����Qgj�H	����΄���E�a9��0���6d��im���pQ�|:N��_G�+A��Nf��eX++�{��UU��$��#��:~���|{�t`��) ��3gL��+g�N�y���w�w�ٌzp�K���.�2���"x��<�\33ֶ��T=Ր݋�!�:\���U��r��n�W�8�2�makg��lܟҒ����E��w��I��!�� �| !%�t8K�j$**��F��X�%I�vWm�x��I2���Ōv�C�	Gf�����=L��y#H��$�=d��QVWfvtC�싷u��)�C�G�9���z8�xW8���_a��*����Ly��J�������lÉؐ���$�\�-�6��^��dw7��n�^_��#���|��Ç7ت�:��42�3�Y<�
����i�(���>6����Vo�R`�����v���}�g����zg6����=��2=���g6��ҟ��iw��H�y�o�n%�Ú��D�U�~�m �����A��vIɞ������$�GF�ރ��(Q�{p��Y� ���F���D9��:�����S�0|F!cc�mv���i��c�R�ݿ�
�G+	�wZL�J}"0ߦ�5L�Gu�}J�����ۛ���ҵ&W��?(�$:٨@��VM>��b'��'\>\�w=��|F����<�1�#e�E�p;��y��;퐊Ƅx~}�o�;�E�F���#˅f2&�_���vw7n;�M$��	��6S f/��jY�\*dZ`缋��t�s�Hc��Z�޶�K��/�ܸB/f�u�p{�*&�����10~M��)���)i���F�4c���@�Ȏ�~o��P�m33�ǧ�����&�i���o��JJ�7?z��V�2��P)���tbJ����	Z&ϭ�g����a������~�V��]8ȵ�zX��uN+�y���[q�ڷM���O����VQ`gVj��o��/-[]N����jkE]ՄQ�0N[�м4:��5Y*go����@�����5��ʙ�I~P����tFF��3f�����Z���H���	�H���:*��_r�:c�͑T���C�>"ȟţȡ� ·�������U55�@uD���ٴ�!�p�D^o�t��^���t���T�Ft1��}0��']��f�x{�w4�v$S�!c�]��iKV��3��7�$�����Xo �ſ�B����hw�W�������������>�Y���j��X_��� ��1Co�Ҝ�E�]�_J�k>��c3�{��\Q#9Eٖ�����z�y�|���Ur��FVV��iʰ����5����������";����	���[���׋r������;�0�(��e�N��y��,ʛ�Mݍ{�u��P�:�GQA� �RQ�"#H�L������t �P̞��� U<nN�l�	�Lw�gS	d�Ȥ���%�����~��zvzW��Nfܗ�e{�����D�������Gr=*>�7^�'\�Q'�����w�Z������e�q���s��kl�	m�+��p��"��2B�c�!�����O����1&�+�:�ݍ/�ѽ������H��x|{�#����3%9�E ES��M��Ƅ66�����a���X���=�K���G�Tb�t��5��P�%XXX ��^����ޣѩ��	8#o�����cc"�D�7�93�]z0��� �_��+������ u�Q��[�[d�1<���%��*=έ�����y����=Bz:���k~�SU�t @L�{�m�}�l��zv Tdm|,f�mf뿼�58���������ҳ������2i��T\\��7LGrB/%B�.�T*�V�k�#sk���"4��7��g�B(>�]���	�|)��"Y<�<�3Yi�B,gYW[����m2Q�56�8a1O:� �ld�sļ�'��t�����xhMPZg��9����u��n����H���K�]lq1ü�x���$g]��|+�c�s�֢����g+�l�W�b�[���hM��#���g��l+鑘�oZ�W���]f�9�����4^��G�	�a��Z~P7���� ��bQ��3�[ӡ�[o����%��\O���?Xl@ۜ,� �~������F�5!��K�rm��+]Q��5�+�.�7�v;S,����DDD��F&&�%o.�����6��L���<����A��^�j� Ł��di��F�ŕ�y�(L!�n�W�#� ۣF������w��_[D�����W������K��-�M�ޟΖ��H��_Y$,&��"��(��-"�LV�ػ{z&�ƕE 6��I>MIK#�N `���^�5.h�o~�,cZ�N�7+�wJp�����|���d�do�|o 0ϸ"'�DD#1:�Jl��F|��=���p���EG>F�@�n�[�J�B(o�I�����X�j$))�޹�!%#˕i������wk`��7
�N�`Y'/7���j��o��Ų��陴a��)��5��Lq;Xl��\^�g�Z�ER�~���[��V�Q;\�ք7�������b\����(�Z�?�ql�(/dK'uW�^kWb�t�eu���\�\Qyލ3���a,�K�v�)���XB��ϯ�f�Q���8}�7P���Ux�2s�f��w3���VD��Xk���&|����q����Z�k}�惱`�����ư04����V_����8�O���w�Y=��cb�j��5Ƒ��-S�h�?+(��/72�Sn.a2�u�ۃ,�6���rd����S����%(0���3xml�{lm:�����|=\Lk~?�ڄ���rm#�1����^1��j�*�N�^G=����tu��>t�hh�B�vu����-��?zKJ�#�h��ׄ����p��0�R��
�Km�y7bj�<7��ʓ�a�I���e�&��T�'�c�� �A�a��XR�z��}S�����U��A� �M@�Z@5��Ww�H	��[Y��R�P�0w�����Sæ	��d�a�@_�`Ʀ�R{�\�ajF�q&k�MB��Y�w�؇-y4��� �����L[��j#�߬��Vh!c��2�����RF��M͍�^�B��*��%�� G��w#�G̭a�9~��cT�м�X�ֲP�ڟl��>c��e�T]���M9ؽ��-����ō�
�i�z�(-]���ǡ��9����p��Úw� k*^Hd�\�OEK x��>lZ]�}���p�LC��L�-��sD|\���k�Zd2q��k���h�ҩ�6�$4����r"�J=$ӑ��f��+1�s�KKJb�m�x�Q�
����|�bb�j�F�v�C��	����/�+���v��A����žZ8�l�{���dޙ{v���C#��;eG���]�a���ˢ����͹��n1��U�ܭ�i�+lW=x����͍�~5x�2��#K�T�}�����K��'9��%��\�^��y����yc� \�/�?6'3-:::"����E��X�v]%����1bX�롾���;O�b�F`_!C��mK+�J�I�	e.̶ ���ә��۔}!S����K�鴯�����06��;1�}:���t'��>��c�pI�uu!�X��٤^:�8�Y��|y����4��P�^����r�ر�j�u7Z?�R�ݮ�5��PY~9���n�	�m�Kj�z� `��F����{s��n��J�:�lU�/j[m��d�ļ~���'Y>��zٗ��6�A'��pp q����㡪|#FC�%���0��c��T*�ȱ�c��3��}�q���ii}\�FF������wAx�,��_+Z�i��������.����
��V���P�����͗L﫿>��~J0�S�-�z�bH^�#�o=�֬��sҐ�]��H:�T�<^�ڙr �n�]ɷY�HָX����Ye��d8_j���U�HpF
n���TX�����l��@��v�l��G{sg��׺�V܇k�A�1��@.(�=S-W��G{�G�-~��B;�C+#s��&�������\ܴZ�O�Ꮚ~���;���e�{�go};�������}}���F�鼏��$�9�����������C�g` ��|���)��P1��|� K^�6��kv66��^��e���W�aꦍ�{�|�Ób��8C�]���*����o����777��Fƨ�#23)j�f��=�%%O�a�F����f(M{���l�=���-������I��B�cb����gq�Y�7Ă�뎣l.\�^���7y���4�ʜ���m�V'��HG� ��~������jA�mR�QNv>qN��P��mW@��TT܃���XT"��[�[R?A< G_���m�>����_����O�'_F�~��&�]�����P�/��vN�q��jc���>C��z/Αυ�~	

�^�\=Q�!5/)h�hK�6%�.�4z	��'''�N��U!�ڿ������B�NW���2-��p�/��Io�6��3��sֶ	��<lt���ϧ]a�2�o�_��j��t� mlw�۱q�'�?��p���[˩����2�Q�H�L�����Ki/K%�bHX�[xX����$�gd�.�(�Y�ϭ���/�^�ш#hu���O�d���M�=�p�*Y�`,QVF=٤����)���w?�|{�j�(���kAR�<?M8���tנoꛘH�ft+Qc+T�$ś����#�.����W*�wr�㬵E/ڢ�í�G|��=��	S힛�k�W��tҔZ������&���?���C�ZU��M;���>屜�����#�n�@L!i�����'��'��W�s�M��,I�_?ЏN����x�!��H��i#�
���8��Y omm��=��8��9��V�Y�׎4qxVJ�ڙ|�(a��E��?�*�Y*�e*Њ�`_@�V����L��z��o���V�����׼G?���)y:���z��Y��m�BWǪޫJ222����	���u	��ttz�
��>���O2� �T���X��y�u�dz��2�~��2�T#멧�b�}�q�.��N����c
/�IR�{��j
��?��|
J�c������t�@�Z�۹��V��w�Ls!x7��=�Vg�g+1g0�b]��Z����GضP�C3?:��aS���^P9*#;#��n�¤U�kD��SYϭ�,�����^��{8��_.����݃��Ϭ�Z�*))}*��*)^�&%@#�QK��U]W���Gh(j\bbv}=������nA11$zz����9޷Wb�*��������?L���ӢB d��L���]�X��wa�t��v���]��[���7���q�S��K%2=!�*�HII��R�����_�s��H��=�tfffx% ?A���ո���nЁ���g6��{J�@���6��7�
G �7�{~��6��~l���-��B�7WȺ�eq�>DL��h#����,Ph���R���j��n|�A-�%ODi�����ܟn��b鳬�^��p����a�v�\��c�<;	�r��}���t����uӢ���� t#�����g$�*�0J}h��J�#����^�
���� ��p=~�QYS�u�ܔ��F�y��^_�OKK{�qf��ŵdO�)�qx4�Q�r�פ�`d��V?�����R��O�����M&���%��YY�3�F՞�qۯ2 ������P�0�������t� �_�ɲ�,���(%���)�ˌs��	$���6��7-�1h�R���S��+���Ғ������H2'���"�|M�.�EG�2#x�:�U&��KmP?���|�BE}�9��y�i��Q^�?[P��rVr��x �� ?��𤆄I���B�H�x��;��c�$V�Uq����ʋ^nn��I��O2��f#�A�Eb�\,`F8k�5�����\�5}�N��.�ʒI�ݩ���"�u����L=���I��M�v��a�?��k����"�l1��>D+���>FD��&��A޳@���u !�"�|pwk�^7/����!�k ��)��M�x�4�9�j�A&끻�g L'��Yj�>����n�����;B��o%�E͗I�ܰo �n�_!�����(^�w�q;�:��oy�3-@�'ጬI�dk�F�L��B[�E[EMM�/��u����#��i��~�9%(�w���dJO5Q��\/��)���g�*.s����B���!�Ǡ�E<x�,��|���f��Ղ�=Q�J�$I�5�Ks`|�"�va����rլ�D�~��6�L���uT3.(8�h�Ñ��:����=�������z��1݆���{�Hz�AR��I�<���LZw�- 0�>s�!)�5D8�� \�
��:�[���u�]���_���F���:�9 Ŋ�:!N&��J��n��q��.<h[z�ys4W�`�q �VB6�EEE����}I,~�)��(��1��8_�c��lOb��/T�`l��R����f�~�������^��5Dn�x�Ba�%y�̓�B�|�]]R~͸g�sz�k��n�nUh�7g�˳��<Ժfj�k��ܱ3+��y
ڱKuZ��_p�6�b���.��߹�&0:�������pk���pYT:������v�C����x$$ג�I-0�ţ��l'm��+��ˍL���1>׃ϕ]5`�IL�Z�!p�Y[[���~hI�kxf��5����S����������qv;��|��%���m;��~Q��pu�r_z<(%%�������X2[����fd\3�pX���#H���5v	�1�.<nO'ݴ��+Ƙ�t�"!��y%r�q�yv�^��̏$"ǚ�����wqA���e��
\�u�cg��~���B�� r�zi�e�����÷�>+g
bϾ|0�UX���3(3$��N�e� Qq��s��0����r�#���o��FN=o��1�hb����}�<�Fv''ރ���\ZI�l&:��~+o��qG�>��A�����G� "����ӗ��N�%s�[I�ג���{@��V���W�v��m8�Ӊ������O�I��{���k&V66�.>>�J�i��4���G)���O+������/�2Eu��/?}.���M���T`�yL��J)1�c����Ҍ�Y���_��v�?�J����ɺ�ي�]�Y_��ɕ0ԥ��b)�ĳJ��)�Y���{�)4a��li�r��[�����(��/ �S�y}�D���'�EjB�z��M<���ͦ�Exmmm���R��'�ܵ���������̧��:;;O5�0Q�)..����8��1u�f�s$�" �G��o��2��B�x�	q��H�����o6J�v���i�����T?��6�Kj�n䤣{��rϿ���v�CD#��{ڠl�����!�(/��>|@)�p�>�7!�@+D��؛C����.,��z<�G�j֕c�p%\'7x�։�����a�i�\��m9�c��C]�_�AЅFllSQQ��[m�Ґ�Xc��n}{�#��L�5S{}Ӽ�zn�(�D)�`&�ݻw9(6�<�;� L���ӥ ��[�� &&&G���sQQ�p�2$t�`�yW፩f��O���}c���Ԯ�Z��=�^#E�uaah�5It4f�
��p+�`g]����3�x��]��j���ED�}����3s��M^я�R	������" �|�����W�Չ�\�<��tu�[��,#������@�`�F�O�R�I�˵D�M���&��,4����J]rTkqi�da���]+fQD1��%/�侠�"���M����RGN�FPzz��3���.�C�����/��.w�T��F�cv�U� �<�����r-������e5ʊB;0+����綵��Y�X��Qo��OG��)�-����춛B��y�ۡ�nZϵA�g���J[άM���2�����˄]��jt�g��=�sYh��B�4����t����]��W~��+u��W�����J�������j�Zk�0�6���%y������ft���rv�{{��}�5��juV�B���`���5t^uOD#`ڌ��ߏۜ��������z�{���2����e� �z�)V�fC��6��`Ft@f�0W*jei	u�2J��q�_��e^I����'��NMOS�YB�(�ʒ�9� ��Z��zw{Ea�7������|��vl2�e��oM�r����P��J��d��c!�7	�`�\�و;Ǘ�ޥ���\���WU��S����7F��R�f���.n6���\����4-�]
��b�
��9$���ol��\���+#�si��&_����E����/10�'+�o�Yx%��?�����q��=����key���P��f���zڀz|�I�gpx�͌p{";P-��ۦU�xx��3���C�rn.��N��+���S�V$P��Y���� ��8\Q�����ۙ�,�����gz�Ԣ�;�Sf<<<(�~ S���ů��y �/̦�	��WW�f�T�^;�
�N"��L��S�J&NkC/�#�C��dvJ�ʁ`�Q��T..��x^��]L��ő���ɫ��͗����u;z���3��gU�IɮMNk�9WX�r��LQ�t���H��c"���������z��hU��-��0��и�+X!�ɢf�ڔ�B[W[+ЊK���ɣ��;�������,d�)�����Ia���Dd] ��,���X�t[?��'qX���C�
������ʕ��jV���g&�-��s���;$%qh���[��A���YMQ�@�"""���~ni��N�&ڎ8]�Ɓ}�y�\��4��>�HM��Y�ח��m�a_���A|���bh5:��!=;�������ݪ.U>��#�Z�Mƞ�.*"����mfv܋�����c�*`#5`��}�u8(����.����a0[o�梥���sbv��\��NƪN�)�Pc6h����E�����P����W�^eһ�R��ʚp�87�MG΢?<�uc��44^�&���õ_�?���(��R��>5�p���LWWT��|ڙ��x�սh�G6|�Vv�����ú��������/!�t�J,�h���,�O�d��ʷo�mZ�4U�=��wޙ�B-�PQV��]�US��ͳ�qs�#C���s��i��ݯ����ʘ��ƛB#�p2ބӟ@�O4�X�����]|?a�7�����GD�r�p7ǋ	��T�4[�vZ$��g$ta�Yk:��Y{Ϡ�� ��� �W�Ť��s��^��uŊ�i|	@�<Ja�oI��79�3�?��_q���X��ҡm@���X	�\���f�nR�<4���hg��&��2�3������E��?;`��L���Vx�r:���'r�{��ƀ���`������Tf#�)��Q_��x����L�t7�������q�/��jw,trR �z������jp�W7�BEB~O.(��U� �(w�T�͋��ڥ��%3�3d���F�*]�y�c�$�M`���ģ��ii.���ǳjC��p����a�7zm�W7�|����mF@P2\�v������?����<��7C$���w�ǪM�|��<1������tc��� qe�W�	*�3B��2��zl�㶍'�`���\|y�ok�{Ǫ�T���'E��o9���mc��q(E:$@d%��Dʡ�\�
cn~��&�'z�22p�A9�Q�G1��&V/O�j��7�QqL�. &���]R�iw�Xv�l�99�j�`_{��P�����!
k>���[����<*�鑄��6�9C���nwR�-�
���PV�.Hk]*���w��>Uڣ���Gݴ�F"�m/� ���[</Y��q��PC��8i1��곎�9ԅ�U�=��z��(���.���!�*����G�o�pf����������w���g��7� 3����*!�@�<�FІ1C5`ή������:��q���Zrr_�D@�kt��&�w⍂�ʀ�D���D�ې�����n4 ��z�Q:�rvvvI|���\|(�Py�����rGH�W�{c���
���k茣?�=�m��8x?�L��}����8�g���u�c�a�}�N��� V郈���n���lo��o�- m��J�++�?f�D������]�<�6sH��%��r�u�x\�J���i�/�Nɩ>P��@:o��J�A}�aE���r昙�̪��	s=%����t'��Σa��7�d;��É�322��X�c�gw߅��Xl�@AB�LP���#`f�7f@H����r��:3s��~�y%t���,.�
��(��aA}�ڄd&gff�x@����~F������ �G���b|�Q��@��������W�555EB:���½���K58ag���Y��ss  oY�H��vv�(
84�g�����	�Gঁ���|k3O
��|���
K2:.�?�p��@Z������U���J���L���55�m��P��j�q�g$ �#&'/���346^�����_C�I����̻��}��CKZ�-�+������f�- ��-Ѷ7�ȭ���?X�)Ĕ�4C��6 3��g�w�D�~�� �z$���7�l��9y�m9[����K��SZZ�k͗�w�i��¨�S��h)��nx& �¢�;�B&���axK����'!�8.)�H�O[��OIig�1��/B/��K��]�!�� �*8��.�ߋ�pފ��S����ƭ\�iV�L,p�fP97=M���g
�z�uķo�/����K����	����4�-^�uͱ7۠@���i}Q[�?B�J��ױ���/^<x��IyI���=v�'99��\%��XZ�Pg���NG&E��NX��c�ji�qq?ۇ�k�6;��Jn��kq~��͆�]��%	��WE�4�8��=����X-D
S_�A<G���ɶ�13cHHH���k[��6�x����iP�A�D$kt=A�0�M�q�l�Ϊdi#d5��Q$&6�T�� _�+�"_�Q ����~�E�V�����^
`bJ^^���y�΋��4R˩�%���!����%��:->��a``x���s�P�_G3�_�K; i.����������0�������	5-+
>P'�m�[�e&�ǟ���D1$�cfeV�,3x�暖6m#O�J��Z��p�6d�\���s�������������}��м�9��8D=�\{��������5�,^c?�wF|�'���KLS�v��[����ɽ¬!���>��5{n(�樗y�Ƃ@,��,���������oO�� B������������G��7��o���?o��W�N���ر�#V�H�Ki,�b�لT�ÇŚ��|�)#��K'(�b�uF����G���q
�Mgn�6�*ʢ�Wȕ���k��������4�s闉� ��=z �>=�%`�|<�7��Z��������v*222��j[���L�1���
=[�����'���JW��
��7�O�u��5}� M�,8�U "�d�v��i�+�(U��Rp�d[��V��ѧ���0��A�iC�]hH��y���p*��R�Y:A�Z4�}>>��Oc4U�<��&]��<i��n��>ю��~�
�ٱ�⮭�c48hY��p�8����k���Y)��u��h5�!-U��ڧ�Ɏ�}�N?=!���SFE�����M�J�+8�"���P�?�o�֛�]���@t"��Dߐ�I���Uվ�z�N�����<7���y���(F�ه>��*O9���q� ͻ-�|����-�<�� *���7|;�ǓX�<==�s��|)��,�pQ�)qС�����;WLr2�K�7���`�2 ��P���6����!��I�9����5���=C�F����7�HC�D�+*����7��$CS�tq�w�+��F�
��m�Y�r�W �Z{\���N�}D�3=q 2�x��� �  ���ɂ:]��`��7b1���-�O���������ttv�d� n2��J�h�|�X5��J$� � �}f� G`^N�+%/U�V����c�������GN�k+4"�������U���"-������lϳ�?4uB�i�|O�J�IH�O��BG+��v�+���-E11JzzT��Q���5����=fr���>�ǳ*eF�mf�\���l�)�>��)}�����t2�����B�5�H<x�а�~h�A�������F`�����%KU�wJJ�Ղ��]��$����%(�v������uvs����,<to�q{�Qf�9���b�ۆ�?K銻��6ɑ�u�����D������P�qiK}��Ow�����]�đ���?��$�a[f䐡��'-5�ֹ^��f����Oqޘptba����aW}�����s%w׾$ᛚz���O���X �lSSS'W�&�����q?'��!".Ui��,��oB̸� yX��(mDFn�N���uϊqz��_���1a]Շ-�wx]�h=������['5-��goi �6I�!�,�����1 WB>�b++-ퟚJ����~�������Ϗ�Y$�������@9��λ��7��P�X���7�;'���xų�ٷq�41f$�$饱��D���l+��'B�fBo�̟��D5e4R������߿{Wߘ��c���4@YQ����c����Y<��f<$�&��a^�us��o>�0���j�<�>X蹠�[K�A
�����@ȁ�g���i�&��/F�K`0߫:1��0�����v�L���3ɵ�=nx�f+F��y��"��γ��e
���b�>�q%ݔr]8U�0�qss# =��	3[2r���=4�*�M�Hd҂zWB�M7��b�e+���+�oee��������1�Wj&�~�c�p�1K�eg\��0]4sQ�Iz�}�}������i�zoجH?n%��*K��&�hp^�ICڥ�����}��<9�9Fg�w�y �c���IRC]in>���|�����jˍ�	�����V�R�oy�3{��3����v�o,���YU���7�&�:7��V{w��s-AIM�CI���s.��>w�L�����]&�b��ֵ�7$��x� ����	===�mb�p����"2�������
��0}狒,Fzz�[��W�mm�r�8�
rjN�}����hj��|��y]�:O���6���I���ëM]M)w�'���\�����eXl43�~>�>��D�������R���@+��(q%�x�;�zN����G"m����uС��
�v\GɁ�h��SY����z	��!D��}Qf��7�vz�����g����e����#c�b�G?z�i��64����.��}���~t|<��;R��`�rg����`|������ *��X�T�h�	�Đ��~�f�� ~웪����Õ�q�t��a�ߠKv���JJEB�={|�Jg�Ʀ.r��!ַ�C������E���b�	�L�|0scN����-�kc��Wkw��L�ydY{)��a����/FFF�:���z��sٯ�^��֢"/��<"6�o@�Cg L:���de�V��{��e��Y���|�������_i�"��ϛ=�<(�j�o�� !� �V��}���as�-_�JU`�.r$${���	5N�@,����,ʜ��R�q�@�WVVV{_��p�\ �h�����!�F��y���Aj��Zn6QB��a��K蟉�»�C�n�2�=�5WOd��]PK�$O5����,����ʒ��� �_��4�ě-ja�j�Y �����m�̖����R��*4Z��+Y���Bۄ>X���_]]A烝p8t��B���y��T��yx$�Fi����5����M����b������a66m��y���*F}"2��͗uTK���l���
]ds��%���PA!X�Q�j8��1EQc���i���b�͡��w<���N6���L�CC/��F�����w�k�V�N�$[��]_�����Ӱ��N�h�|jM��)�h�������ޅ�>�0֌.{?����AMꞈ@�:�y��2������ )�HG�����)2:����TN�;"�̎[c!v}T���S���B�F�7�aƤ�SVRڐ�r��[w�5�~��4f!��j�F��bQ&(/���K!�i��ob"A9�����}�����sК��	����L��tǻ�
���r��7�jUb[������B)M�OX(��jr|��E�/��֨[�p���>̵{E�7^���\���f�8�O�Z��Q���en����C#�+�z�e&] �f�G��d��/P�x_�
�a�A=@J�#�o3��^�[x-�)fM����&�1��Ն�޵�|��wȎ��Ͻ|�;��Nഁ��J_�s�j�P �y�u��>�B�帉�A�$��5QJ����-]:����0|BJF�}�����bxJӅf����g���?~����C�-�����{�ccqnno��	>��a�4Ө�l�aԛ#����Mez+:(��ڽzb�����ܓ�ƅ�`s`�b-��&?U/�C'�_8(]U����^c�C�s�G�T�|�-##C�5p2T��wEQ�x�%�M��J:UoЌ�C�2��#�BBB�CC��|�88~qq���i\TD!a��|Y
�	���"��Z���^nd�,�����_�T�Vym���O��
b&�	e{9�=`\�����5΄oD����9=����*�`�G��X_�0�Fħ'��,:�233w����"!�0U�+��&~A=�7�VCCQ���_}ڧ'�F�|g"��M���������n�0�Vu~��ͶN��D��C���'�r�����x�A����"W��Ą�5�b�>�w�$$$`9_�?�#��qZ���;t������Ӝ%(HO�q�j������IZ@F�=�>���Nz��*���A�J�X�z@�}L5t؝f�v$J�/Q�j�p�@���p��}(�̊HGG���t����Nb�������̼���?=}Gi˔�FC(�d��H�X���5�JJ}�.^���x��
���^�o�{G�*U�����&���?����y�k^�KK���������F6� Jˬ�����8� DReޏ��*?q��d�x&�4R��.�P�^���G		�'�w7%***�/�����7���=��S/�H��$�~����wG~pr���`a����K���W����ǖ�Y��<xĶ��ط�ح����Gn���r+�ŋ"厎������Q��Dxx��M @^�c+T� �h��h������t��h�)����H��pv?cn���r��/@ǹ2��c���9��	Z'S���4��?��}; #u�������#��r-�����Q�8��Y@�J��}�K��`�Vg��M��<tk+�/��k�e�E�n����S�������y�/V��� $E�䜳��Sa�&���cl��"��ݺ���a-޷�W63U,� ?4AP}�S���E�@`��f��読�&�L#�����(��vv���=�>%��h7�1go��A�����*��P ��<�q�z���`�U:+V�E��¡�+���b�0�A���Y��FYVV�7�'���Յӥ�[[�_�ġ�Wڤ�)qq����4
2�ns��6���T<w`�;^L w������3�=�R�����q����9��FR�~���n��p���μ��د�W��"�K�.���$�x�n���E��f��z��|z��b ���0D���rp�w�'������	03Gٽ��E���L\���)�`1���V�|����f���� d��B�6��'
�R���a6�s�����ڟT��c[�(�n=V?�@8533�Ŧ�-Ȳ]�����Bd~Y��1=������ϱ�?
���9~
��KG�x{Z�{\�pck5H��xa2�u�P��o?z��|���#HLX:ώ��Ix���N���_��⾕�_�8��G))���W2_`���8����.N'Xlѧ�t�d��_��2}��d��mVv߷8,�忿t�+�5~��y��!�����>�z)>���{GǷ�wW ��f,�@{�FW��&-r��wv�Hg���p�5.U����<�-��Rޝ�����߿QP�'���n;;�~.���S��g$da�'~�{~�]b���
�樰�t��AD�.����L�#TY����=����T-�����>��ٸ��ql-���#�q|e� ���GV+���&v��|�+���������?�3^�����ط@��_HHh����_�m��Y�:��%3��Oy�c�ۄ�`�_�����a�>�x��90p6�K��;�[T|VY��*����ԁ�Qo>���\k:� ������Ӓg��H�(�u������6�5Mq͓>M���MK�����Ж�#4ٌ�'84�ʌ)^��섃�ap��z]52"���'H+X��60�,ۘ.h�>����������/�ъ��Z����� ��|	鮪QA��Ѹ͵���ې�wc���Zx�I���ȫ��D�L���¯��Ӱv��5A�WNd��>d����_���ǚ�@�~���A�2V��G̟x������鹸���� �X����/6:�N����c�#�QCR�t'��.����*�I�>��ᕘ��
W��C������Q�ƺi-�H��+7�_�/{�cj������H`r=	B��Z��\������v�����#����M`��X��@�7f#/ML�����wv��+�x�Z�p��*�WlfI�m�,dj���^�O}��v�Ґ��2�����:=���A���Y%%��!CC�D���"��EqhXK�V�_�����i5��q>�G��?��2,��kQ�AQB��n���n����n���������o���~����g֜1�f-��>�]���3��B�����?^���u�i�t]\|�O����
� ^F***)u��0{��<��Kևۚ��׶�������%%#�+�?  ��� ������$��O���dK��D�TF�~9�diSrHkw����_x�`�逈�(a3Ֆ�P%<����i6F����o��
�#�\ȯ��VY��!{b�����s�%��x>̀Cau��4.�������,tj�g=1���P^��6�c١Җ0�@��~�N
uN��s��t Sy����؁ƢS�����}�`lLS�h�= p�������y�����&��
.\(������ۃs��q6k�=py��on��% � ��Y���c� � �^ٺfz�,_�Xg78d�I��5:z�p��؟��q�6rd������������ЪT�#%]3�O�8@BFft{p:Vl���|ԣ��������L0.�m~� V26�����e�K�^,�}�q�`gJa/�uK6��{�w�ܑ8�<����I@g5�I��d���mYS���S�ࡃ,��,,Z���D����w]]�O8(�oצ�lq�9�('
Ր#E|$ٵ�ml0��ʬN7�!����+����� ��U+�I�|����;���� �r������J�D���:����U{`�hI�=9xƂܳ�&�l���O</��׻��º\��(����V�7&��׮
G�b^e#5U�������� BkS�HH�CIm`���Q����`*++�����9�x��B%�r��f^	lV_����:�W�B�T��mNj�\��:�!���7>�z��\�3���	ʝ/���J��F㹘�5@�i����u���t{�&/��;���9��(�$N�21���Z��V��s||�^�gX���]��C�B�7���j��ȥ݉��t����Ƀ�7���y8f��������y|�l*��p� xdt��vO1_�b'��ݷG��Zt45���e9PP��s�W��
�ZJ�ԡ���ֶ�<`=��z�ա0=����an(��5U�iDxx����,�DŮd�㈊�[�WW����bn�o��)(>�Ȅy��O���x�Sx�wBC5���P*Ro4��˻c&jjj�l�m�	85�8_[��E)nP01ax=Gm��ǚ�¼u8U{����qb"����`��d���J�Z��Ǧ�s�\&��c?+��ä[p�$�keɟ+I��̓��.}�'��dQ/.��S���;��a>8�TPo��7��r�g�DR+hO�+�b�#d�C���Q�Z��� �U\�Z���&���ׯ5ZA���	��=x�jWHhbb��c%�S����͵�~�t��2=A�$�&&�&�r?��������N����ˡ�W l�\��_1H[�r:��"��=�^ UD,0��Ҳ&����7��B󪲲�q>��x�ii�z_A���l5ʀrm�w��,�2%{�����&,�{M���v�[2��w{�Ϸ������x~����S`�(*Z"�}�1aoecQ^Y5�(u����j��Ie/�BrDZ.C���P��"_��!H��z>u�tzj@�/I�08�iR/� tҠ�R��j�:�o��q�Qm,L�[C�0��޵���P�r�2ֻ����`�siB�6�X]]]�����E��a|�e��,���g@eI76D����a�/}||J�����|�6�M�
���9g��H�h]���Od;7�ם�:_k�ʩ���V���3�\����,݆�0a�]�=;[�Y.����˽�O���NGs�}�{z��������p��{�"-a�T�%��²�BZM��rWݒ�Х?ҥW�{��p�H��EaM�|�I�"�����~g��Sgλa���8��{��{1���\*���H)��u.��m'D{�g�Jǩf���Ċ5[`{���)*z���-�m��G������ [�N�����¿��!���߿Gy�h�k$��]#?.�%���3v����Ĥ������00���$�,|��Ϳ.��:�Omm��1�֓K����r��b����s���7�:�SNI·��V���Z����YlQQRB�a)�J�\��+*(/��r^�W����^�`bh3��_]̫���dg7wa3:_�C[)�f;�Ͼ�������2n�fr�畧Dx-���?����������H�EMd2�$_��Z!�8�MMᠡ�Et�l��= H����A�ن[]�DI��Ȁ�qb4�I�]���C�(�o+����n��s_Q���h��p�8^���ø.0k�vv�No��ɧ7_��X�a����VSK��L恊��Oʩ�V�0�Q���aC�@�EE�B��@�K��ǳ�'<<<�i���6���@$�'M@�{i�{��mTFE����!F0����e��ʳ
�^g���31����j��t�(��uA~.>���İn����^�蝣Y��Μ�V����ڦ?�a?�������������ю����bb�veI0K��˼%�/���_Z���UU������[[���ʸ�r��iii}q*<�A�<�	u�u�w����r%y��������� ��:Q�R�pJD���"�Č?}n0թ�d��(�1PW�M���l'''P�̀�i�����l�Z[y�������Յ��%q9�B�@@di�(�C<Yq}�I�ť�o��o����??>�SV033�	�u�Q��QoK���K�Mmդ`D���Z�]E&���?��x^O�����W����]m=�ٜ��텉���22�����-��6ܮ�V?-Q�d+Y���pp�b�7<��1�͖\�8Z禾X-6�_����㭗���������[Z�7:���S���;�M<כ�ʬ�Y���yb��� ��藋X�S�7j�d�WHX���{����7}��Z��HXAp��R�`5/���/��Q����ֆ����*"�)|~�ٓ���ǚ��iB��)�m&����Ңе��' ҭkl�WF���"L+�5x����\pA�
`^�ֶ6 ]�{���枙"	՝�m<����s��GK�>����)#'�QJV���]�Sn����Z����!���ΰ�}bbJ]��es��q�>>>�p��<�TPP��^SU�"�	��/�]m�̸����zzu�Ϧ�҉!���-�ӱ'����ٹ�\ez�XN�����SS��.н'�F9�נT�dn��9n��ă
�II�
a�p�v�(�z�������b�tq1M0de�#�̑�P$T���ԽE*B9UcE����9�&��$��gh�������:1!����@ypڻO�`s���k�zj�̅����7e���y޿s?��pg+���	���о��&$&�Ľd�k��l��M�Q��%��$�*���8�~dfdKd�}6�W��4�!����e���[�*hrrr=�����r�P7e�K���h�}S��m����>����wt�1�PW������'�<�"�0�%.n`s���5�06��%�8<���=�!��qhhh�,T��@����80�j���7����x��~�Wג�,b\�||\n�L�����3`���|��N��	�6���q�<���I0��0�*L�X�� �������`����չL�Z�!��8x���NT"ְ��%�C��r��p�k���N�t�"""�6-��������^3b&��M��ND}�T�xxZi)S�C�|2��gY��� �?9��`�e,����wu�*���_��⨊56rdfN��A|�ꕇ����KJQQ�p8��m8)��1+��![:��6��/�O���P���d`������S�0�����L�<��2.���p�f�W�v��.���N<�4j,�'.iVsl>WWn���x=�6\�(&6���#�pSN���mC����usD�ј��gK�\�b�����]sv�~a�ɻΪ�O����\8ߝ�u~@-Pa�8pLA��rg �B�;h�[�MI�ZU�6;�^2}�a�?�/___��'��s�.���U��[y�A����P�^���o_�w$�]�����kllQK�����:b!!�f�t���A����8�M�>ջ��FѼd� sYbKk7o�.X����|��#5�xkgG�𱗾	���!�'���5�%����p�r�?+�6�?�z��[�GF9�������P<B���99������ �D�D��d����������/*�}%b��L�ߑL"z�TU��}�H|�x�B�j��۷���p�-��é���?��Ưcjk١"� D�9�Ɓz6v�nc�l�POi�a[{{{+j�������`���v�ȈLKmj�t�E�d6����x���	%��T�?׸���Xm��<�'�6(g���,:�f�LVÂ���+Z).�cd�f��Pý�&^m��P�'�]&X��,����<�4�o�Ya�݅��0�d�j13�C����$���&�m�䴯��5\O	vV,�=���-<����/�g*^��^���JJ��ƕ�0fJ&��g��s�����Y�yL�{x���QA��zZHHH�$z�󧇮py<�?y6��9`ˌ�������{��i7oE��.�N�Bd�p�E>�蜘��ǔ-�V�Wߓ�Z�p@��6ICP�\��}�|��~ST����껠 :L�0�^9��	��gf:�e�$Ms�Sio��F珓8����) �^^O׏�>��*��ݪ[+�ee|߾A0�,�
�N��
ADb�[��������S ��>.���q@��*�j-�|4{+���6V8yrzJYEb�]���j��dQmb����M�W	�h��?+%������zw���⢜L~�lX@]>!�]��BB��BN����>�)&F���no�(��^h�ڈ5]��o�=��Z�6i��f㆛zt_m�Ea������*���A�~�T��:zɛ,���3� ��A���А{-;�5mJJ
�N<hd���8�WBQ��	 ��6�dd¦C�J9;?��F�jYb��⛜�����iĬ���VN�y���ji�����rC����zJ⫸����L�ع�1=NG��*�]�͡:7����� �I��G�e�w�r��~�P�}� L�L�����(�j�G?SR����*��w�ܻ��W�Nb����tU��C:�g52:z@q��\�*�8<������/\���0����?��Zm/00<�$��������Ng��*n����7��r�]e�H��M���\�|���ۻ^������ᴔ���*��_�$GEuV� 3��'N���T����Ư�����XVVV��|Z��������<��_�>OMK�I�11�����bw��X��z9g�����k��
��N�_��^��B@FF����,�/:��k,,�^�|���U�p����|�|��������v������4��Z�ڰ Z�A=4�#���giɔq�l{(�)''gc��-w�#X^�DTTH��o�HK��=��%����0}GP�4F$!!)V��&'G�ʊ���jK_�t)�w0R�
��Sh�����h	�	v�A�ۗ!I�_v�m&g��H��%̵"�4����Ҩ�'��TV�$Uc8	.��ܜy��]?���9�:ֱ�>o3�����_g�.T�[Z_���ZX��f'���q�p]�!�v�oZ_<M�7��0;�\/n���Я!����'�*#�t�fomD���X�g'Z,d�%Iu��C@m!�>����Ƴ��u+���������clllqi�Jmf^^�ʊ��N�"M_���C�u���sj��f`����sЛ`,����]`!+�Â���2�f�Xˑ���NV��)�l�d8���՝�C�PU5���C`6��z`{
�z�:���|�3�%Px.�C������I3rr���Ѷ�EP���ƥC��M�1�]�]s`�	TtA7�wDC��s��d0�P1!�n�EFF�b�#3�����)Վ�P^���!�΁FQ��-*�����@崹F�X3���8�3�0�8!CC�rI�=6k]�9�/C��Ʃ	���$$�6�t��w�W����yǲ�PA��Fڇ�?�sb�C$���(������2vH*)����La(P����ئ��yƥ��1;��F�05�]�`4A��3���2��d�a���iA(((W��]���v}����444/�����Y��ZY�&P�.�O���h}�#��*���fW�-�s���_4�@�5��[�/..��,��נ�����J�r�]��)@��H���EJ�Yz��M����I~-�K�M�_ed0
��23���}�����I�N�
uy���s�0���s�.6��c�:ցw
.N7�*㎯���o����j(�jp�G?�#G��:�Ij���v�y��(FS��l��09	$D�V�G����11�9/�X�c�(���A3�qKf�iR��"��pל��O3���EDN��5���������,������ ��m���"6�:�b㜟R�Qg٭�L�X,��5�t�p$ǋ������d�� ٮ�P\Un�����*n�@� 3<<|�-�%%��Sբ��f�I��P���$tt�f�qA�Oh?��LBF� �C~i):!7���G�á��Wn/��b�����; �F2�#  �;���H�U݁A�Hh��6K��TU�\�7s�8&!6?������~@���ﯯ�!M����>V�_̀��JtE����QQe�5�3j?[l�\�{A�x�cH%��#��j��_�o�n�'�}�q/W�Z9H�C2�`���l�
��0��|�����z�;H�-$Kf�W�&���������:�|ʊ�TC �Ә�+/5��Kr�}�����5V$�1����ͮ���0���;���~A]��]p�A$�8QQQc�������	�{���  ��U3N��2�.����П.}��it�m��������h}z���"|y�;����ɯ������А���J���Duڰ��y�����r'�r��	�t�е�6��WJ��L���h�r����H5�݇�˶�@�jjk�����գef�NNN���-�"��{{{/pp�~ �^�N�y��9*��?^.�uj
��ё������9�M������L�N�+���tggg�¬�tM�.�����vv����_v�;��|� ��VI@�C�9	w@�/�������B)�`�����>���f�5e�Phc�����t�撺�k$���r�_!2-�},�a�v}��w�Ɩ�T[]a�S"���2��HT�T��L<��H��B<�,�/---�H��_������k3n��&��ѝ�PO��p�K����v�+��������������9_��<E�����L\��vV�_?���
#xBBB�;r�cH+�L�8\��}��� Q[\^�V{�>��V��ui����P�A ]�]n��/����3�Af �J��t{�R���[��o/� >�ON� �H�P�K�更�a(�bk��z���G�+�[��U888NV���{�(�3�:ێ���|�c��X32�N��ۋ}d������ćI7(�������U������ �ܯ��zg�a����3_k�9�j2����ws㋰0"�D|�G{�ɀqő�z�k�CN��Ni��78����4�Ǎ ��z�z�7�3��"�?�H���d`a����^��"}����V$�����M�ն�H�VY@I�p�B����qY��c8��T���n����
2،S/��iV;�M�~� g�BKL��Fi��C�1��w))iJ����ǈ"�:�H}�h0���Y�`�k`ѭ)���srs�.1H��&:Q�%�d�<OV"�U���������y|<�\��jC,	���ʀy�_���p/]� �����eL�C�<D.����{���צ��CؠqW��)��W�U�䜜o���Wk;�K�
�8f���^�8��o �]};\hX����>��\\$���Q�~��yX����|G.�i|���ņ�Ӆq��
C��}R<~t]���?8x��8����=Q�瑱˙c�v4?23���0!�r��\��q��p�)sr(�D��$8:���*mW9nǒ��-��ҁ-_J��l���^$)�yt1�J��0ǅ�`|���6�t�'ه	�QdX��uſ�Gš<ϙ�_WW�/�~�r������tۻmY�E����i����n Q�������#?�}�����keu]���*w���T��$3�'B�ܘ����I�}Ȁ�K��1�����j��ɬpx&JJDz�����и��ծ��~�n�#�E(�l�bjJQ�խ��xE ���L8��7j22�U�r��$���h����:A�x�����֙ [%{�����)�r��WW�lF=Z4�UF�q���G�ICC#��]"A�c�"�L�)�����<��|%�_�o��Yì~<��v���Ѹ:��;��7�L`#9�?��^筫�G��c�|2�x͗^�,xY��u��B��6�y�Ⳬ�Zv�s��ضU�8J~����p)iJ��s ��9 ��z��~n�;����s��I�Uj.���()W1bds��5��QQ��/w'�6������&n\�ߍ�	�|mCZ�hkc���������X�����D�>)�1�H8��b�q?�_j s���p_��p}�~�����g3�1��|6����ZYs�3�k������'%7I2��(�����6O���+M�{./E���A�_v����x5�i��`�̔[k�sr��S`g띒C��Q,��X�?5�7b����;��%�nx06��W�1D���zҏ�ڸ_D�_���j4NT�p����������b�8^���K&��W0S����<��}^0�~9>���Q�-�"�hF�����W��`�
6��&`��:Yp�A�{��S��S�%"�G���y���kl�Q� QQQc�;۲�($:gq���222�_�2T��l̅󀺬��,6%���i��H�����4��x���|u�9sy}�4�%I�dtwҌ\ @�аub����f �jF��$��9SS��+TXt~v�ifF?�����G������	����\m���K*����e�V7R��jw._qvc)x�F���l�4�T��0@��"<=�67�T9B��cDZ��o�SoU҄���m.\����?2j���%��:�N����pֈ7�x�<��y!���߸p˘��������Z�:��򣤤�j��w����kk�

7����1s�N �̴$�@��4�b�,"�_h�����''����A��A�S������F$=���9�t�fu� ��Ap	�c�va���؟%y�*��!��� �������k��J�˃_/I�qf���{���W�S�ܻ�M.>��(//��p�K��ɝ,�Kх8p�2�n	�0�����:���6t]ŀ� �c�j&�.77�oL��^�H�eB���կ��k�^O�+̸]2'�2���"/]I�h��+��l˄��J�.��6Z�j�52�>CDAI�Y	���l.c-�����f��Ų��ֹ+��de�����LP,hrt;fF�ة9}��/�<����N��ױ�����U@Ev@�ހu��̨�\��T�hN�7*�>�N���{��\��~Kݍ0�XXX��+>�ѼB����a�D�Ю�IE��C��ߏho�HFFGWk:���B��+���W2k� ���H�߾��ёy��!v4���gg�ZZ<l5�w͏f����tLL��m~� ��H���p<p׈%��ڹr�a���`����}���D�c�Yc�io�Bt���z}�"UY1@CJ]���@�u�O�|�N9@a[2��1a�ZfC�~)���&v*�uLO�<�ꒁѐ;@5#�>���`d¢�|��?�/V���2��gF!ф��7��QL�Ԡ��x?.��+��H��-��l����N�
2-I�G��o.ƻ�0бU5���m��v�� V`:�� Ī1s��vL"{�ꝒB4XLbhWoo�j�ɘ���-�Vn`��/
 ��c�VP Ų�,���䲀'>��	YUUu(C{jz:�d����4�C-�5Rψ��F�G	����t���a������?������s탹gVǣ6M�b�^,����Y����Ճ�rDdƭ�{.ք�M�}�q����*^�2��^��^�:y�#�l�Nt��~�A��ƥ�.Hj���N����gõ���'���d�C=�s��U�� �D*�����il��l�s|s�eu�!���SiP]�n�_�kcx��ߊ߾!�E�\.���V"�VU�\�LHL8��0�������_k&����n'Do�#'���n�d�~��uQVV�e{���D*K����B�E�GZ��˙J�  6��㄄�~s����ߝ��?>pA� $Z����z�k�NIb�������\k�˒����寍&3Ƴd�$px��V]$�����+ŵ+)ǔ�k5]��SV|����X�ç��B �2:R�ݚ�g3VЅ�9 4m�sVh~�p���Tt��;))�7H���9h����S����x�^�R�:�e�-j�XQ��lU����Tԥr��:�@�\
����ꌜԲ��]������c����5���ID��n�ʐE.�M)(����h �ë{��jk�$�.5U��4SL\�Jբ+���_�缼��E�%�c9��@��@%�{����9��]������ize��@��4�vc*��/�h-��V���+�=��������ܥ����	��(/�W�U儂���f�/�%���“��t/*-	y늴*�UYSQ=�PQ�9��	��������R�ǻW�J�%�;]�	o�����ɤ���'�"�

���ϢI�ճ0 �p��`�[��"�cH�XTQ�dBrX1�����A�������b$����f�\"�(�7~|�c�S�?�o#���)vvv���G�_3��K��~�24���AEAUL����46F!''�6.`�wQ�?}xx���j퉤~_�i�?�T8XG+��66�I�.�gg�suv����B�����U,AaTq���1q����k�.��@iC���,�bA��Y�]+ U�F2�L��v_���jl:3��s�M���';�BA\T6q�$q���۔�r��}�m�T���4�Z���	�����d,8F������Ǐ�%DF�47������u��#���{�������j������R�\���.�NAM=2�[ .-<����r�׶~t���o��Zr����t_X��Z��Sr�����|hXi�Rh@4	��y�4����@���ixx�q���2��C��K	�;�+�ޟ?�M�\��#���"--e"�k��"#��c�����5�����\�[0`������&9���S�D!�TT����|�lZ%z�@A��)�S�ueu�J��ma��}i������v������׾?������t���+��;S__�70O�hbz��6�3��� C1c�!Vlj66�չ��c~�Wb�!2�͹~��_庨~,0e��Տ�W�]�&U.��3x�X���,��o�)I�>y2w��� O���K��e�fg��O/\�%4���d��
R�jtz]N����p�H���^1o�LO4^+	�T>m��͹:�X�B��ܮ22"b��PY��b�u<S<��򡧶�O>Λ7�`�޵?�5�B␮�C��{�{���4���������/�?گ���@��h����bcqyy;0:�?�̆d��;���HY����CgA�Ä��TMR�'nb7˧��������U@ ������|��EEV���9yl	�yk>�$���`3�@7��z���PsswB'�:����«,6�b��G}Mg���ñf���򪈏#�'�x�ܰ�R����Y9T�nnnN�WbB�0����w�3O�@��-4�l�W�_���1>E�����ǟV�(q���L�ۅ�~Y+��ıO��Q04|�/_�7?�t��s��&_�`w�PƉB����p��ё�N���f�x��R��5��"��Pvz�Q�a$Ԑ �����C=ᯰ0� �))�J����������*o`qN8�萔�S�fq{pN����	ی#������n�����r�a��dKKK������;9����,d�58>66 3q����+`d�Aԧ�ָ޳K$s��A'���H�|��U���H�������B������#�6�\ww�c�I�����?�nH|Ih���|D!6Lѳl���I./N���s���/_�����Ϛ�ދ��������E��c�2U"G��C�'��c�mĥ���<��1\Li�Z.j�-Uc�[:���5�gӃ���}}�*J����^�~�i�Y�:�[��H��|Sa��Q�[�:��Л���\�w`�3����������dn^T$>�'��"�� 	���@��nԐ�������j��L�]c�[iE�虖[�&޾�#�$0�nv�)����Nn?���j���Z������A����)L3�ܣ�s#燻7���Վ�;�|P���|8d�?��	�ɮ�7�Ʋ����N�i��ʚ�3��x���zu�8&���`v���ɪ1QV铒�����j��񆄓kq��� K����xl���������i���~�Po4�`����D��7���C�3'?����2-���+@�X[R?I")��!au�1�Z�Ϩ��L�u��\ý9�7�"pMZ���P6���`[�Ȱ��	�pF_@�BfR�DD)-�dO.}W׺�U5�,�Οoʻ�OOW�,��J&.H�/.6��.�������[M����K���)|~#�i����Kꪪ���3��>�����(�������>��N�����������:#`���-�T`5o.�����'���8تo`��琞��]�؝I�I`J��xn0S��<:�keBjj�u�}������?%��x������+EN���`|e��8�3q�K6�);R�V�۫�!���RR�e��H���,,,��U��m?���%�.l�.��H�8�(����?g)c������z0G�l�����i�.󍦙#����߾�3?ն]�8D999���/gj���������vH�_(e�މ�^�:*K�oj���l�����%Q�W�۴�͚p�����vq񘬬��Ϊ`Is�5YYZ��7���$%��t�_[ATE��U�P,L#��ۯe���\?�j�$%-���s�ف��v�zj��l��B8hE�}�Р�����J;b!Kmm�'�5���c�<��1ma!�w�m�B}�.|a�3�0Ƨㅘӆ�?�04"#khd��p�Xj�YN���,��fϴĪ�=�����JCS�x���bu�o��#ageA���]���]���F'/��R�0UB��+2��JJ��;.�V	u���R��?*L�g�K�ޘ.�����:���[�Ѷi-7~�R�D�W��L�0�,�w"����j:���0.==��F�+U\�f�%�În�t���ϯ�\������������Wj333}���E���������{<�ǵV~/̀�������(*�0}��`K�T������5b���:��P�8�388i�F�7o��7&  "�I�ϝ�ܜ�T�ڛ�] ��vR	�^Y�"���ag����;��d�?��e�v��0��ja�@�5	O %ҊAгI�� ���|����{jbw{	�1Oq������#"�̭��I�
e	��!���<y�T�;29*�;4ax����:O�bI�Z��c[o�d��A���Gש�Ra,�c��h�uh�K���!�X�*�^�Sx4�2~O���#������}�E�A�.7�)�t�D�{�r
���ULv��7���9���+�3�:m�<*�����6�T}�������j8�AM(��j������zǛ.%�~��mnNu��4p{���tǿ��x�u�37SʹzD
�=  QFF���ܰ� �����b�k{GG˟�������E�\#yR�����W��Y�K柮��I�����A���k4������S'�ƅA��&Ӂ�Ǆ�� �\�7 �?::�lhH5hz���ܷ̀�m	t�̌	�����¦Wv:O5,��j�^�@�/gg����ͫu���6�d�f���x���b@U��.�a�����Ku���V)=폵9Ҙ����������^��#��*�I�,���#��CB�o�0�mW5���N��=X>��p�ɷ���{^MI��l���q�*Td�=����~ؘY0
��WR�y��{���WQ!-/6]�����ƛ͖)��B�>}­KM���O�8GS�o�{^����x�l�嚐���,I�84E��F�7o��������+}w�U$��z��a��q7��i���Y��`?��ӜҲ<:���{�C{kk��Gpy��d��F���WWIBK^C�>�w�=��PJY�����d{�'ᱱ��~
� ��ZM����0��es�ЎPF>�3b����1� ��N��^Yq(����@u�����,?����6��:J� KB+�Y�YAiLo�f�F�u �{�-������W�v����L��m���htLV͎�l�Q��0��.4��7:��CMnnI��߿�:���KJ������B[c
E�-��k�ss	yPc�Z��;���=U2Ξ@|���$����0��T�����a������=@���Q򘸸T��`g����&B �^]i�RPd�z���[mwH`ii�")�:v�r2���� �e��UT��	8�4S���_N��L|cVT*��cr �?Y��*���@���f�.=^��E�	����y
q�o�F�'��\?�w�}�rX>�����!�|���>Sa$�W'uh�F!��E�3$j�ź%�H8��)����CL�ƻ���6����1�0=,H��W��.�E��i���勳�k���&�.^���A�A����1��J�䔬�z��4T�����R�xrt�̒�,2������܏B�:���+�~u��t�j��������a��l�e��~ 26�Qz�NqU�_CCC3#��쑟Oc@W������ӧ% �2C���s���; X�����&�MJ
��I\NP�y��*�~L���h���r�鰼����!�o�<n�s5VP�`��Xꥅ+���$�����W������ �Oi����T 766��}���z��h"�urh(��G��@2O��0M(9�%T�AV[G�%�d�JDD��i�0�W˃��ڵu���Q23l�a�biC,J+3��l�M�e��	^$ ��ّ��F�S��˛��۽�&�r��,c����Y��w�"��8Y���&�KK�)ǭM�;���x�J�Dd�����9�b�|.B���A�zx�B"��wN��Rϣ���g�˗���:���x_a}�U�T����~���my/�����&+k[SM������N\��Y%:&3���'^��|D�d�z�*Ҽe����)��yO���������x#*�������i������$����w��ah�ܳQCV�lg<�٬�W~�gP;
 ���0;-E��"(((�].��� ̀�v��������a�����:�ageņnɁ@�,�6�[P@`��zC�X��	f��p-���G+�?߲apss�z�.�4�r�?�����֖�L<�{���tm�������6�lll�Tt��$����SĲrr?�UXLg'�m+�3���ρ�m��j������N?.�<�!,�v��q����U%e8
�^�U��+C@�[|y���v2j	����P���Ŷ�a�敼eL&�o\]]�o�V�fI`�H�<E�Q��^���%�U|aw7m5�xQ~ncaZ���9	��Y���WJ�ϞQ�a�J]m��Z�����u~e�
|���W�u�b���dD�:�]�Ǝ~o���]�����Yx�I��u8�mt��NLLT���Y�&q,ڿK�s�(���͒"�ggg�����2=I���N$�?ʎ϶e�-�B���?QQo���U3rrq�6�æ��)a���� �Ylm午�"��WQ���P) F�g� ��Yyo�bŠ��m}ޝ(Hɻm
���谿��*��7�����x88�mmO��(@�����˕v8}����[tECC�:E9^�!��ͅ�����T^�Q��h��k�X12 $]:t��� �c��;AS&+Lf+�O�v���2��>��U����(�xo�����ӳ3k���8>>J���
%��}����7���%��Ϝ�?��׿��h@�c��UmtV��o���tR22�D��T�Z�!;A �T��?�r���:R&����2�TD�w47w1���c�����
�����[BG��D�o�ux[F�x�[[��Tw���.�4�Hq
��l�zf����	u��X���a �TrδT\4���������S�Q���&p�s�$�5���}tu32�	y���];�Ǿx�l�(�?�khg�p�����zf�c�����]M*oQn�ɀf3
�WYL�(����X��ܔ��L��C�AL�k��b��7k���W vO�HV��J�BAI�r!&��_!EQcN��Vdx��XV3�}1Dr��+�5P�~���}���CACq)�@��XJ�������F__�������799 a�8+���汃��*+;9�vh�ԡcT�621��J�q��Q7�R�6��Iyi�J*:ZJڼ��E�=�

MKcc��0�TT=�r���۹M���w����ĉ"��>�Yq&h(e����y��ǿ���K*��5e�o��/�����d�e�K�t� ˣ|r� �H���z6�)րR�T�$p���+'����J�&�+/~�����CE@�l��K}g&�&ܬ:a0XN35����`y�5�����O�f|B����j��s��W�^9�_��P��=:��w����쬽�����V8t �DE����(EJ6/�����������i�^���%twweE[:*����,��3��?t��K��|����ᢆ���
���sz��3����G)�
�V�Ng[i�!����LN*���� ./��
���utd�@��,���"rr���V�.zO�w��E���0��YEE!��������Ś�0ш�
?1_q9��jr��F��g�L׼͒L^:8PO��G}�XM������ [ �
\P3ٙ����*vI]n�A����d�U�_��s�*�g��:��V~qJR���eUx�9��lȢj��jM�+�P�ń�z��N���?��*�f�)��	�����	)�.A�����nAZ�F:��C�;���{���9k�.����{?�3�goz$h�����G�L`�KKK�_d�N�q:E�=�.̦҇U��7��v,�5$�.Qj�M�Ԕ~�`~��+��-{�F���h�<{���u{䪔]<w\YߞE��"���6�E��0��aE���J#?�������7�̇��v�	��0� Nj��"���.��|�8R*�i�ff~��.			�S���� z�QTR�Ǧ�(��^g�]肷�R�<YK�x?�t���k�o��!ddd0�]���_3	�ʂ�Y(��;K®[J��]ln�v�l�|���ws��z�O2'DE�a2��W���p���Ɖ?�8Mc��^���	�Ω"��d�f�����k���{��-}#5���a�:�3*�<� Yx���:M�/(,<���8Y�J|����N�`7v���
_6�{Yuvb!��?��+�*���AQTv	�d�O��^i;����>�&�VWWo�p/�{�:��oW��a5 ������c�pr��RK��k6{@!=_��W�m�{�rzJ떊q"��9�]�}!�@����D�~�laa��4�Ç�i/�0M��6נӼw=����ru�7�
)�������˭Gf~�|�j5�b��D`�u�~�Sx�?��򨧣foN���|1+�8~dn��Hxp�������z�V���7y����!��A����X�E�I+�i��S!(H��9�%���������e���TTX �]��+ �͋]C4h7k�o?�m�$ǁ�����C0Ҽ�FFڀ� [d��!���M�� ��#�u���V��TUU��������>�Q`�^�_�/)�D��h���o
����xi�Rgw� щ�
5��VxH��������~&��1,<�ac��l@9v�H�62������n�9��Ѻ5�cw@wVF�n�E'���[d��E
bol�h���O`�л`;��W��߿
K�p�rg)��ڼ�*�����^։ݷ�+Ǧ�xRD�����v�B�)(*Q8X�?��ϼ���nbn�X��/1��Q'X�/���C�<*.9�!�=�q0�� ��\�0���LD���|� ��������q���`����o<Ӧxj��/��.��#�ԭ���|�+�v��h{e�� 3M�Җ~�v#ىvs���%���U0��d/���ȸ?�~{w7��'י�.a�f~�F�y�����Ʋ��+�V��*��B?�+s��&���xz���H�:����p���Y�*;,�AP�Ĳ�%V.�@`�@���p]���N{ս>^��r�I�>9l9��B<�էF�!����A��#��v7	�i�s5����7 ���������T����q?�N(O�g��~�L|~q-�˨xbTL����c�"����:�%+�o�(
l���	J�/��d(eS��~���=z�{d>`�`Y��QO�W����Y`P�FJJ*���rq�������]Y��t�ڹy?]����Ժpkr�/��&d�ga	v2��k0h��)Aqss�><�8�u��U����\x��q�ÙU?mmC���J�;__E�>y��R0���r	��ii��I&&&���������S*�b�ֵ�����洙ng�<wYM�0c��r���jz��a�
��_�~Ů����Ӄ,���H�t(	�H�=�EW�i���os�����"��{,��ϷĈ��>��v���|55�x��m �V�ad�4K)� ��uʟ�u�y99�a���G��OK��Q��L�[��6��N�1�ժ���s�>~k��0�o�
����O{�!����b�.:R���װ=z:���]	��}鲔�J��5Gv-���9���B��>"�Q5�W�~��U��@*�^�o444X]f�،��0'GBqB��8A@҄$��"�1<I�т�L��!T@����bbT��3tm���YY����,J~�nX> ���&j%?o#�2+t�w��y��Q�"�yVn.�R�:>�;:�v� xuC)��.���>�k7�����ip$�� Iv�2�ı��aO�V��N��z���c-ii���taa���rx
��<Gf���E�Ӱ������'t��'WJ��vH�����'��CSaSk ��;l�^�v12X-B�"��T�5��`sy``!�fa|����$#m��#Z����<_���KL[:�zg_8Q��+A�K� ��w#88JTVVV)?X�1�դ��#d�΀��ƁBf��c$ߍ�����W�ݞ,[���NU�k8]����������be�����*q@<��x����qΗ�����{/������2��6�m{�:NMM����"O t100���������{���>�pߜ�����|��ڔ�`D~wM}�$���ܕ��tX]K`�� `
�ի/���?kkkk"��,�/�}\:��9�ya���U+F&��w�P�E����v��zw�pU(AO���C�[DO���^��+S����i����179��ǎ)Vsɶfo�� �%R�W��қq�5���c��4p��?T�Xz2�K��{P7�Y���Oַ�La��yxP�����D;}�� |`vf�{}�U_cam��񨔸1_���c�AϚ۳.�.�����Ր�O	K�9�n�t�����UWĞ��d����Q��2����+ߎ�f	���<i����)���Ϡ ��w	5,Ǧ'������l�J�V/-��f�g�N_{ܛ�PS�گ8XK�ukW%��K��7t�Z~H�I[8�sAj��]Ǘ���5�mMШ�$<*�������,����8܈�5ӂK����TUE;��A0���7��!-#���w'�~k}u�PE-���) �����z�����_z������vɈ�x��Z{��@N�Hq�����M�AA�ev�T���X�m[��}h��;���y�4��-��'����
��R�������`O�Lj[~;
�f��D�Y��GD�
BK>x���}]����ƳoE�
zpE�^��#��A��+��:��ҫ��~�k����6Dwឋ��Թ�owG,�x���555���V�nX9!L
o�n����-S�%�F���:�C]EB�~p��}�ѣ؃�k�U2�d�:.MKɣ���T�>���Z@v��q�{���|X��`�ソ"��_����w���zmdW���#f(6������hs��E���}Ѱ ��*�1;�[������>��G=���Ҳ��2dN��&f��~�G�}WF
�FrlHQ���/ĺ�n��U�i�HUW7�y�Uv���P����pDCu���K�NRve;�G���0�qS���?I.���5�rvq�z@O�� C��Ű�Ӥ�?��ce�W2Ղcc�2��B�{lj��jn��w�K�q���}Cٲg����̬,X�ޞ�J"o�N�y�t�ұ�+nX3��l��&/Ogݖ��N����� ٞa����O��C��s�"c$`�i<�0+��2���M�a9���6k`d�7��y!����� n3Q�������?,�W
��3�3�m1�C�R2>WA����!�A�Q&��R��0	�=�yd����U(	��{K�����@!~�P-�``�b&�x�n}�{ߠ���淔�M3^i7�,��G\�@/�{��N�Z����`�Q���T�-+.A~U�{�jFR�T�>�R=vs֓��`+C�TO�,,���:j�AF�:�z���Y �f���՝܀}�B��<����)����}�ۙo\�׊�25�V���5z�ѓ�g����Q������l�����J����Y"�ř�.X:��G��R�����;^3	��	e`���ۇ�6�g13	��Χ���v糧�f����{�u#������Wx�a��+������������8GnsG��m_܏��/��>��D?\��4��F崌�c��&2��m��f}�3)S�+(�Nʗ��)�P�x��۔��Ҽ��%� G��$!�d��D%�(����7�CX<<<���lzO�c�L����������$�K7�Nk1<��I�Y^��Uذ�~]�A�H���i6m�鐊�?��]��v_�܃�>�0�����|��4��9�An�#j#�}�����o��]?���\R����MWSa��nD�^����5����/��f
:�����ms^;�~X��H +; 4Mz����#EE��E�7(L̦�t��N������wz��m;!�saa�7"3����*F,*A��5T	��m�#�7�S~
Z�*���os������i��M�
��ʵ����=��k�p=�5��Wht���Ƶ#���0���}�Yǂ#��Y�;CD���D�j�^`^�K��SA�����;H҉�Ͼ��>��KG�M��׫\��f��H�Z���`O[�;##ø3�E��[�*�B��廵kP�q�u����� �
�9 )�~�0�6��v�~+�xĜ��Wc��2ݎ������L�Զ���v:���
�FT�5rwA��i;]f p����®W��.9|�A�á�������E��˫gK�&'��aXe�"���rM �

:۴��w�j�5�i�^������u��,Q[]�ԁO-�@꺨z�]6�v���ʩ�jx(�#��͸CS��$ ��i��3���?�*�v	����%		d�㤰�:Sƞ��PdҼ=yw�_FB�e�Yll����}�-��ű�Η�M����z4�D�ț��s`e8��s��cSSi�f���&#//1�}�t����5	�"�!V��&���U��f�²1^�+̰�,��<H��50"�1_N����X�<��秨y���a�Fe|��mA�Jr��A��Q���7��dbm�+����Q�m��G<�AS�j��������ho��ay��6�?;bNv��^�H��#^�M�s�:���>��B9[h�zi��O�j�o��pMD*e��V+�?��T�Zf|5&m�l@D��YrE6�3� �P���0=;��x��\�ݴ�F��E�FF��vL���wR�ñ{ao3�� l�s��� ���l�l�P�:��Y�&����a�Tk���!%e�l+�HGϊ��i��K�������E(��ˏ����� �+Os/��e��"㗽\Y�Iw5.��|/ب,�B�w��������Y~�-�Ϛ��#�Ǐ�� N���w9%���s<����%ia�����71��Ӽ�Ia��>��ehh�]e}�m��ݜ�K�����Ի��}u#�Q$�v�F'*J\��ヰKII��VV^��������C�7��[�98��D�h�3?�:=}�� ��!,�;?oT,�g���v��&�����~�Ug5��������1��ٹ�)�L}ɀ2zd~��06��܇����㣘�^)ٗ�F� ~���.��ֳ���=910�G����]�W`�*	B���ϮSYp��G��<I�t���H!����Ω���˪W�'��D�s��	H�	j�FZb�3Wj�v���Ɛ`yP T�S��Trw</���c�OrۿYa7�9Y��H�>�vbo�[[��"�G�jGi.���$s��U�����&I4�ͼv7d��
��:��S #�B'￞$in�x�E�Z���E���]L��"gkFMa�a�/����ZF��#kU�� l����~�����u�L_F�	"S@� �.4­ֿ�U�����n<"��Kx�Cc�)�ߝEG�s���"��{�l_79���L�"i��w����b�揗8Dя^o9s�0�Z\�-��íi�߿�	9fL���U��t�@��}�	��J�ٷ)����(����#$y斖�@ޚεÔ��|�@�?�IzK?h}�>��\g��>k\�wG�����C�p�Q�p���̅s��O�'�Ό�:2��(�jk�uLD���E�j{w�����M��s21�)�%�02nɭ�exu�qA�]�,�˄�++k�_j��R���j9Qo�|l{~)�Z�Oh���H��*��}�?�+0�UN{QV�P�a���K8.�+�D]Lظ��<�ʲX�͟��	�ވâ��uCc��z��D<9D����Ʃ��DBd�8�.���s��~���$��>�pt|�l�gl����y �B/�Y�I��wL���~5���j���l�<.�0�]i++V�Z�)�ɞ3`�ɋk:!��Ԅ���MQ�Tl��S����-]��=n�V,�:�t�HS_����i6����q����hj~\2�;11�_��̷����ut+lr*����w��z�����6�:A}���[�0���Kt|�m���� �A��e�����v���{	|�o����IZn�W���8=ڊ���5}��}�������ё����w�>^���8���!�r��>8$'''..�#�y��5��x^^^��7M�̸M�Pl&??̳�ť�����*��߯���UT���!njJ��kC �Z�dxx�?����k��4��+�eT�(77�YkX#�w:�`E3�N�9�E��~R�K�7�������̴G3�ΚIII�b�B����,���3�'�|k8�MB#���/�� ���M��ڕ~k?:%���Epp�h��D��?��ehH3�����ڈ����hok+W�<�-+�Հd�|��N�����-�4{�x�Y�`-���H�EViqqD�/`L~��~�"HUF�_v;ٖ'kzS���H����999�ddd� ���<�⺷8fDNY�����-���~��I��_vj�x���ޑz!�S&���t�AW[�;S{�jW.i��lξ5��۲�|�lR �Δ�6�z��LJ��u#���k����Y��<�ggg�`�=988c��4�z���
��[�'5�H@��'@�i�Ar�(�^�7jjnn6~�Ћaoϯ���������j��;�Ro�=)�W��,C�R��S~ Z�`��rA�����s(�`1�X�̾E�����S�[��a���g�݅��3��:j0�{��˱\� ,e<4�9`"���do)(��o@ ����<a肧��53�e� � ���WRV�
8,�&�����J����ׯ�JI�&eBw�쳬4X�!��8�&;O��o`�-VXS#�Q)9$G=(�eߩZ|�X�P_?��ٓ\`��4Pa!7��rrr�|�NN��?'��*\��k^��*��WrY��2���r~�k(����fK� ~���V�������	&�F��f76½�׌����x.#mm2IIɨ��G�T��k�6f��B����{-�(͒H�vy��.�y���tQJwlkW���C� +��i������yMII	�����:�����,6�
�gc�I����) +����vfe%�s 8��鍋e���)�q4����E�w-�3����	���cbf6<r�m	!5,n9v=����D�Ly�Zg��{|g�ܜ���(9�'ß~4o~�꺶1V�h-�!���\�^,�R{���������g	������^���]aq*�g��bn<�RA�(3CEE��_BSS3��Ql|����wi*��H�By�oll��� ]�vMPD�g<��]�z@�@Ժ�����;��>$��T1���#�����>�	�xT����i�;��>���ؔ���W�?�\3b���/�S[�n�H��LIB�g��̜x�����619)�5dM@NlWw�����k��C;V�=3l|�� �b������j]���8�|��/��*[�����D�gE���E�7�[�ȏ��#�7k����4v�_����i�A���x,�a�i:էDB�ӭ��C^a;�IKKx�R��i[���~���Z�Y���|K�;�ڡ�\2�۹�m�����s���ؚ{�E�@h�d��˗�����'�[��a�-Nح��L�2����=��(��� v_}�O�W�����bm��z�,[H���}v ���rJu�����꺜y�vU��D�'%l��u�{����(�g�F�|�mx�r ޙ���6�h7�����F���=���� �jnxy�r�@���������X��������QlP�@1I�9׻�>��,���&Tx<�.0L|r+���g������a�������,\�[�J*���z��I���߾������8^2�q�����r偵���� �;=���*:ff٬G��>}���Q�7���@�����SI�UU|yyy,a����P�K�@V��~��#�ݻw��ߖօ��z��-<��u	����4�'��DD(��~N 0����FR��M=br��+枝�V��"_�EV1C4��Z��z�b���^�uA\bb�YCI�ͯ���h`�s����P������3��YYz3b�MM��rx$/�ofC��=X����!�$��W�3��c�.����**�����^z<H�� ���WM���'�b�^�VbJ�P��L�.���0��/]6��F�m� ������R	��0��S]s�	��dPCB�~>"�W���;"������Y�[��!�&{!���t޻��.O��⭈O��4�_��T@��!2��'an���� �5*t�t�=a!�t��8�M�����/SS��l�?�SRE�DP��º�#����:m�S��r�p����Y�&I��T�F�	��b�:��)�t�Z�#'at"�>@K,��-l�V�p ������2� ��wu�0Wkp���s��b����,�"! �]��r;��622���N$:&&T|1�^m\�w H���J*e:>zu�C8��G����~���7?C����^,����֝,R"�Q諴3���bbb1���5�8 �`�`Y�����
�oZ ��<�ڱb���8>=�������.,�rqq��N�>�\洍�j�|�
[�*XH_�`v~��pg�3F�1��u��#{T��(��X�|&�,�� ��i�UZ@�7��4��>�996o2qr�DGG���..�!���o��(�':��-,��RA��� y�ch_��So���+ � �����pE����,�d �J� �{ �yxx �8�� Q`�����Ŭ��?G��5}j���g�	t$%�	`�C!�8��Z�g@ck������w�XXmo˄S4�->��I@�ԗN��
��"���o�����+��/���ɉ*�[.`��p<�р7��v?evy֥�W��Y����"U����N�(R��>�WH��d���5��b��Ǹ�U���}V��9���#j<�����@g������ ���2-*)��=V�!:<<���\D�@<zD��"��Q6����7I��s�C�2[��L'��[[�__�l����p:��ly�F��}�`�+h��]�/,�F�����u�e��Z�_�f�@�+�;;���Y1�(�5��ݏ��ݑ/���i�dmo���#���0k�k����g-�������}����9P�SVZNpl���tll]�Ϝ7'�'?�����Ӑ�	}��`��*�_����1:mv�Iz��_?�gT�K3i��F��u(���z�����)/�tf���;w�<�,V�r���,$"��FG��²�S���#�$$|vX'"� ğjW�5LM��~�o����Ŝ���
wPa{��b��1��e6? '��������* �M@�NMM)S1ܹCe=��H?�L�����.�7n��v/{���ќe�qC�J[:��d�sf��}��F�&�.����\𭧇��PAA!�����I�G�TYY�������A �Aw���G"�vs�;{ݷ����[��e�� ��[��zb��]N����k^g;����j[1��N��$�BQN����Z����Ym��M x�p�A�d�s�ׯ��k�����,�	�$�N�`P��� �0�r5y���O��I�r���U'��,���>9���|$�2��'''�5�\pW!#�Q[Gv(�=��Dz74�]��-��Nh�%�x}�
񁴤��7obhJ��� �p�hŨ�,��ԡ ��L
�aJkJ�b�Ak����,����B1��@q��)?Da��c`RA�ᗖl��dpe�ーb�����[�Ch�ۜ�l|������R ���R��lXc:���q!(�����0ܾ]:VDd�;��ZBb���ns{o���R.喭 ���S�8֛D��f�r4������ �ڝ(�ˑ�>������(�;Ŭ??L�X���}���>��x�B��D��F_�ktM�����_�K��4G,
���@*�2���2:`� � eN!$$�C��F�ȈF��2��O �����}Ļ�M(�Yqz��~�ސ���Û (HQP\���[S��KP�í���1۫y�i���AW���q� �r���а�����=��I�Q�r���]\<ڣ�C]`�%��6%��n�+'gk�thXw�6�����+�Ȓ�94�4����oa'jד�s �`( P9D�>Z���̢jhh��i�}\>y�^������$�q�Z|9����5�>>H�\0���z$�a�Vgg�o}�wy���D5ܥ�����چP$�����b�P]
DU<vvs�]}�b3����A�	��'�]��sZ �W�7�_�z��N$Sv��2܎��<�"O.�T�~:^��o���}����MSo�̆�-X �˿)+(ܓ���3srr�2R��&x��g}~~~=�� �O ���d �(8��pO7<S��6���?�܆mu��
j>�$���>�()�w���}+�2c�oU. �3ɵ&��)��(?�8|��1+���5<CZ�º��
�ٳ}d�,�=�>{�� ���� �rZZ�j-?7���	&&f�GwS���<�#���#���pJfI��,s���/�mt�V�Ѱ��\A�i��{�>��*b�lZe�,TW�M��ݘ�'�`wo�/E9G��J�{��r�&&�d򙘬�<����5�djaw,8��X���D�*��]�m�<,j��{�⮮9J#�(=D�>1��N����� ��N�?~��[�������y͍�`��T*2���\QL�H0ٹTn=O�F�Y���j��>m�@-�;0)]�o��Y�YyT�CZ܏�ɒ�Q�w��s����!0^ރ��A[l�u/�ƃ\�Oj9*jji.|q�������YȈ�G�M�6�=�wd��� ,�1s���m�XT��������:�7�>�׌r+���sʬ�a��|��|�~=�*���:X�PꙙF�m���`����=k2[�f4�'obf�ׯ�a(�6��e�g�9��!�-]��g�Mi�R��ױN����9aŔ8NzM��${[�U4$� �4�и�S�ѥ~a����ZE�u�H�RK�$|m��F�bb�7F睿X�}�~�S���2�Q�J�h�R��%~� 6��)�@7�:��j倗=�"����.��w��-o���i�Q.�
�`bd|"J�����jˊ�M�H��&������M�5n��r��*
�1#c�7��m�@��Q�<[���Z�Xj�q�&�W�3hWZ�8x����1t`�k�|I��c��2O�����M�m[[N�e��2�U�J57�~��)\�p�&,"���ٌ���|~yW�����\���n�-�#}�}�3�Ѩ�&��t5�:1`��E����H>`WU�'�Z�	UX�>K1�ʏ{�?��+]J'�3�gw��� �,,�����k��,n	��r�}tP97�//&ځ�B�R��h�f� /
m����9P��u��JB(����!ܻo�/�f������S
��g*�QO�Y��D� o\��B	���~��8%`iM�,� e���qp�����6�թ�a��Q�>��S^��[wF�46�888f��Ы�#jL��e��ͦ�|�EAG���Y�N(r�x�N����囍�'����,!�<ѩ��3n��6-pu�|7�.���nd8��再��x򈞮�e�Y@f��ggg=����Ԯ�hw���K�*--mޙo�][cs"�s�}��OD�
����.��C�ԟqd�ГۄK6�/y�����HC�޹�uR�;�B��G��h$~����wIFy��T^U'C4�lB#�߾��k+�`Q뺗Km��9db��1�a}~a�c�-ɸ�?�`s�<�N�k�W"�?���ݿ:������JV*L�i�0y�3�Ⱦ�n��o,�����dnPq�����-�i �_d�`�X�Ї�.�[X�嶿��*�c@��^���P�n|�8[��g�.�A��*�rX�ʚ�	ԫ�����"���b����}X��j9����/��.�mN���S���ȥ�
'&'��/kT ���1 i,��'Ht��|�/пw9��R�O��o4��G $QY��8ݲ���_Ͳ���Đ�lJ�^׼�BF/C���������;��ϖpR����j_�ь`�S�9�}q��P�dS9WM��P��/���[�cd���(0����j�ۚ���xZ�q����o�@���]��a�&9�W���,W�]����U�i<� �I�Y�9���n̾(��uB�_��c�'�y��ɠ����l@vmЁ�+������E~:>{�;���^L�p~g~~�z���+@�՗�ۻ�z�(�1`����~ 6��3f<[�866�>�}��f�
�W�P�>��w8Y�Ie��g)�qR�-)����P�ֺ��`�����0,��ߡ�B�[f|M]�n�	���Ǽ@!��;7���L�o��0޳�3�����\Gåѷ ����͙��o��p�흝M3�~ܞ��n���z�ۭ�v���?�wt�������Ex">,֛�e�
�� ���1�#	E�T�5X��NH�v���f������:�{xKk+������x�׈{]�A��TT��ENM�G}��	��{
�n�����ݢ1�x"�_�M���5� �������$ۿc�4f7�3qm��^^���T��+r��t �����1��K�2�U�H���]Zsm��]>�X埞��ծ"\ɮ�I�s��%B�+�Q�}�-�u������f�����9��1��FR��o��N<��ï��s�4�?�������yG���B.�T���-Ρ{�����_�ON������Q������^(MOg ��p�����D��<�xqS�U�B��wY��#X�䳸���S�+>��#b���)�m�0��B�W+����쥾'�_ihm��������!,�s=��@�|:"�r'ori�D�{n�٥���`�X{c;A:�Az=���'��;X�����3
	�U�z���{�'�	;�����f�>qt5���5BA რ#��C�ќ	`5`+��o#)C�>�/���j����$J�YҋU�0��X(XT����|�1{�m4�T��!� ���=��i�d:��O�����o���4_,)-�LLT�&++��Jp�-��1k��:$͒r�[����>z�
�Q�h:���! [����~SM�XW�r�yMr���so��� 	ɧD9���^��/G0��&&�Q�\`�i�0�.m�aQ1����qc��̵`�����i�� ,�ǣ��dpO����	Q�F�W���Y�?yJ�E��l��P�2F�0��*����N>ҡ>1[���lu�Zv�Q$c �E䬂$.�D����K��~5/�� 

���x����g� �c�E��^11i�eI�߈,i8�;CG'����׆��*��ž�a�T23W\I�w��L����<�ɖq
2a�*׽��2�b2���3�	"����3%��9�q`�����`������A$����
�g �����c��d|\��aS�g�MCY Y�|++�1<����4��脢槈��q.�s2�8I�0��Ç��S)X�a��X�IF;��<B>�d�`�����1�-0|�c��&�t;'�y�.�:sJN!B҆W`� 7�m�%���;���[��W _>��A-�^�fY]���#��4�C��u����T3_�d{��M1#1#����W����^U�k��sAo��CV␐(x��PQW�>h��ce���'�Yq��� �Zݛ�f8xx@����o	:oR�� ��F���0V!��{H6ڦ�5�o��>���чp	dcN�M_�x&�5�k�<l\u��o8X���2\�g°�3�R�rW����R׾�>n��pR���^�$�����MAZM��u��ň�3P�R�8�-;ߵ�<Q%���^�K��|�ܪu�ݓ1���P������)�����j��'�J�&��U$��3�PL���^��377�a|xG�r�}v��6���]oܨ5�� ��`����nЁ��t��CC���ԥ�gk�U�c_u.����I7k�sE\Ӹ�q���hdlY�nahDD@8N���7����$�����<�������V�\NZ`V?���!uNKź��~����ߢ�&ЃH"B	����LDR̴�D̠��� �������~�Q6"��h!�N{��k*�ޭ�#��Y�\�b��ˋ��ъk���6
�_�{� �Y�\��L�#���_v :���44��.V��7�i��_A�E��0e�aFx�ޜ��t+�����E���4���I#�B�uu)&&&Z"$�r>�JIa� ���uB9U,��=�r*�᫾H�3?tө�*A-�»%G������9� ���C��oPC4����>����s����p�]�w��@U�xt�0x���2"�4|�O���# =}�>V/MC�/"|3���z�a��-�c+��͜(>v�g�M�0��iX���n���'��,f�͉���WrmiiT�s�|VU]��e6V��3��D���s����h�n�y��i������_ƧO�6���e���"���u�ٙ��<7��EZ�C��܇*�����H��@$QF��9�^^��l�@��~���$��N
�������Q�v�Ѧ��mާcD�k������!�Lɘ�"}DD�G�0�2_O ��D��jLن9�@B���I0�����d/?��F���j1Kt�+>��I6�M�x>[H��Ԝ�H��: o��W�5��rHӝ&j����^
�VT��A�ہϾw?�|�R�}�U{��gU/��/�]��/s��˻�A�D��5�����>�L��֤<g��8m}߻��`_����8���T�B@�a�(TC��?_]��|�u�NE� Ϭ�CE�^���\�\D�i��瞧����ظ8�A|8n����D�{���D�$�:�
��*�W쾵�&~C}�/������A���k1L�k�+�(��f)�+��}��&>(��J��#\�_M��0������7��@��` ߐg�������j���������F�X� j	����K��z��Z}l��&�M��{N&Wu3�NV3��/�� 66�)�M
R��cE��\�3�R������b>E"�i��Y4�����*����:��"f���P�(�ow�G(a�Zޯ��������d=�N���]C�G�2�	����󕢁�T/'2G��1:��>��A�8���iFt��7�!N���U]d���HTH�UG��s4��_u'��D�(��Q{ 9nږ�VDG�/��]ÛqĦm�����w�>�j>@��%G�qFx���5�~5)�� x:0��G
;�.;��4,��X.����������2���8��b�����j�,đ���^Z�r��*\|a�b���'��#����A�;<H�^ؒ��)J�T��f唖�o���K�1Mv�t��\fZ8��b������S�;s��)�9k��*i��5Z�����p�<h�0Yu��,|�1�c���_̈��ˮ�ζ���d�e���A�4*9���j�����yRU��xb���69�?iB�/�@M��?o��Ҩ��݃�T��/����8X8�JJJ�#bRS���1pqiq����O�|xf>Ɍo��V�F���k�oH��Ӗݍ/�����')�k��w���`<��T�i�/��I��	#����9(6g7��;["$�+���w,������[N��'}�e"�^@�f/*Q��y ��G��|�҈']A$�X�a��׾�g�#�GJ��AW~��������_C
�uC�9_�d�<�&�kyK��5���r�#1�g`<̶�9�=i�/�"ΰ��N�+H�H��g��x��)��մ�@>
RE�f���Iw���lON��7�����Lz�+w�'r��'�i�"D�	ں�5����v
o��Q�^�͢*fHȋ�ۺ�c�j�A�xe���@�'�����oP��P7��hK@OD&{\˾ȼ�y3T�ddT��V
�x9�{����%ߣ�ߝ	h�����֠��}
��C�N]}Vl�j�
R�����|�o���q��~X����,,��|�I���;�Y�p��Z��MUy�-�[��g��/���j����d��R �5$\�������3}Z��:F�� ���+G�r���<=> ^�`2�p��hc��ѝ*9n0�[�VQ��i���m1%�j�!��PCNC���^��n�Q��Y�3�Q�gT�_By��}���BZ�I������|��X�ү$?�:n�*Ϲ�E�Îa�J��J�-A8.�R�w ]��]r)��]6�l_�l�:42� �Јj�#Q�GHh6x�6*I��M%����z�ч�o{E�O靨�|�|٥^�H{�����j�(�4����>y�4�pp_?[9���֣��zN��9�&�n(��:���%�*|r"O:�ښ�V�r�Ȗ��~��RuNNN�Z���G��'}M�{yK����t��C���������̸D��Ь2��=��"9RpVS��'�B���@�����"!n{(����a�͜r[!��p=��w=�l�������B���^LF
(�VJ��x4��Xs-���n\$�����:�"k�n�쵣znwKK!eN����3�Z�)��e�/G��Z�����ǌ�Կ,�Z*Y� ��Zt��)��tu��b�B��������#�0JLd ������<�?;0���D��r���Tҡ������845&���^�Of{�'ˀ::li�Pc@��ã��bY�!�m���������F������-�i��-��M���{u�\H�J��㬒�\�}�)=})�������X�0���(�VP�zPL�b�[���/�~��23��m��~G,�<t� �����5�
���"��o�PH������mi���.��YZ�a����|M�D�8A��'$zi'k�qbꑂ#������Y<`l�j�oF�s�<��z�D���t=�\�i�Y���)�e�����CA�G_�-��:pK˭l�s����z���]��L���������B(>R�9C?=z�p1/X>S��uR�WSC����c%Ԋ�D�����}��-:Tu�1���["Lq��^����5}i��YE��f�ܹ�,V��`���(��ݧud�G�A�~�ⶶ��_��(����4�]
�7�֒�������Ӻ��f�v`�5�Og7����\�S���ɦ�8�+$��I9S�����B5@@��M��i|kik��`��s���+����&��c����'�R�S�,dw�d�H������7{�蜠Q��47PqG'kW�Y�ϣ��N�1����9.w�5mFSg�k#�{8�ni��z{"n����l��3K��o�>�u�gKM�����e!ٜ�Sp�5� |'�D�5�+���,��Đ"oE��w�KX��;:�UQ��n�� ��B�|U���j����;ѳ�}5��f	%��FJhٺU��܊_>�d��x7�^8#�b#�ɷ���a5Y\��ü�;�N��k�]�G��C�W�E���.,����HI�K������4H)��)   ݠ��K/("�t,�t/H7�,~��q��}�93��[��;s��\Yl�,,m�Ǵ��p�d�"Z���Tw��5��cN�£U�S���RЄ��������]���*�>�M��L����}P~	ս���<貫����kz��������k���Es� t٭yeO`�cv3xiCʄ�a$(�j��hN783�Q��Ŝ�v�\��>c�wp��[�2M8Uff&�_,\���2��Y4$�豍�P��#�T3�s��`2���M��Y�Iv�׎<�R����<�d^�w65H�?XJn�Tl� ��^+ǁ����o��7ȓ�0�G	�iA:��A���V~^^^����?}�T=M�CWt{kk��	������;/X\H�B��&�<�:ՠF?�'K��M�I��=suy��'�"l�D�Ġ]Gϸ�r6mRz�U��J�KF��ҙs�G�E��v�y9�q�4��8c͙��u�9�gS�}�Ϟ��O&ǚ]͒#��x������u h6\m���"a4�t�<�_3r��c���%��-��Q����am��/KM��ɡEY�$����|44�IEttt\Y)�jы7��Z��H��z1��m���0{�q���LG�o��KNs�,�cFn���͠dc��u7(E���`����������<Qg�f�t%���]2���� ��'	
�@^?H_���p��&�:��ڡ�Y}�Z�+��Uqn���|�q<�ݶ�'m<⅋xU>�A�&
�]x��h�T��I��Nʓ�G��q(mOڕ	�! D���J��\[��Lcݪ���4G��p��ר�ro���&%��|87�Nd�JP��#4��l���ł�(W�X ��b,>ˬC�4oJ���ר,>�!��x�K��S!f�ޝ/�t��7A�H����gY,����l�A��Ţ�)4z��f}�)��l9%C^���R8�W�@���ߍ����S��h�p�+c`BeUU�ZR!��s�`���H!�A(���)�TmH��Ŷ���J�Ƒ�����ӱ��vZSFEѨ�m������ճ��6E�D�:�t���%]���6��Y|ߢn��r	i �r�� w�3���Ԕ���Є]Y���7�G�0=cwj��pH��A��('�^��/�~��g<���L�k榗�Ɉ�7)�3cGME6k�+�;��}��̂���7q�U�<>�=2c*WK������-D��d�^�ͱH�q�'��	���ܬ5��r����������,���KO�:b֓��~L��a5�?[��,���q7R�0�����,�
]�<��cK��@'��q`�KP05
��f�v/�F�9���3ʕ8�[��s��
I������� ��,�Di�p�:����h�략YJo���8I�����;w�|&��Lx�{b����?<J�w���B�����&YG��lՅ(i�T�B3��D���î��;�tf��x�8B3�eH���74���-�Oڙ�yد��S�ؗ�^�;�9O9�pߩ	A�R@�(K?�:#�U�A�E��>�)<�0�/r���3��D;( O���2�8è�E�.l�U虉	��N� �|��E������$s��A`�#X�+q�bP�!N,u�*"yH����y��P-U�ꤟ���ZF�Yt���x'�	/���� ���:d�WB�|4Y9��Ч(逼?�}����g����1�'F�\�Qk�[ƥ��s��v�HZ!�?9J�y^f�G��S�m�a���{�U���?�:.�j4���N��]x�)�ocn���]�l�*S�����"��W�\���eyc�L�L'j��X<o��;qé{v~g4l��,Z�>Bv��o��+�iӭc4��Ê�7�A�q��B�ft�Q�{s
���r���,s�����������7mΘrl����y�^���_[[��R�ָ�J��fE�h�[��PK�����x�e�<���T)mC�Yg�7$C�RkV>kc��àB��2N��N�-�X����ů��W$��%��}����`�f}�丕��k{~�X�Z��O&E@����&q*�Wި3��Vt�ф]W@��>���/��O9n_dūp�p���޸�LUu�\__ʔ��A�i	��d�e3��S�'b~�3�f���O H��|�m1��0k��ꈗDQ4U���-�;����J���C']Z��aO" L�r�Ը�TG�f��z�L@
��ܪ�8
��NmJ��B)�M;����&%�x��h7�W���dʵ�7����2���	� �󕎾�.�K)�n��I��55����H$woy�f�Zè%�+���初�Ĉga����8�H���M��;�x���E��=ΦsUH� ��~eZe�����D��II�}��_.7���\�!ӷש�
�-$�66�����i���|}=�Ӓ��\ ~� T ��X��b�ʧ�Mm8ᐾ�+�8t���U���Y[�m6��Q��V3b����s�NJh^��Qp���	/IY8I�Sq�]��⿘r�H�>ϱ������B����m-  `Y5�Դᠭ�2������x�a�^���1��[���Y���q��=?N��*�����Ʋ��8�r0H�l�|�����@i�*ݍ���o�|
i�/.P��_Q�W��Fm�V�˱y_שu���Fho�ܭh�x�̷ҽ w��<��\���ڭ��z4�����Қ�w��k������c�q��_)�[]TS�e[{�5����V]��l�TKOO�5������mC���G&����f?�60b�W�%~1Y����6�ʶ(�<���)ϕ��f��7,G �lN%�.�d������<j��%��p�4�!>����iJ=��×���W�3�]��/���D��j4��P�3���p}h�o�x���|�u����js�"��dmtxxxcV�n�j-�/_�;|���� �B����7��������s;��$�T5���_i�/7��뽺�{Y=�"���5��~Z��`NJ�>K����e�]�s�~8�� =��~Pt����L��K�WU;=��	����P�BUj@�ƋCd3�ތ���3�p� %a9���kХH[ƿ�vI��x�m����E��b`�K^�����5�>�r���O�+�%O��M�����"B_9��OE�wu.��/��W���z������NyQ�^ߏ��W)�]���Z�Y�;I4H�Et藻v6`�+�N�I����ȚY���-�x�x1Ag�f���i���+��|J�~/.�<��-��'���F 9h���	R��S~�Eͬ�}���|�w���ϊ<Ts��U��8�?nL�f�������9���6�+̂`� h�b��=��Z��IU��� �l�1l�g^".��� 2�L���;����M�@Fnҹ�H�@��d�+�A5�����欐�K�G�b�;����t�#D�qܰ��b{�˾��u�+f����b��c{�䃂�qy��.�{c�=$:�C�}�$m^x��q�v�(���#c�EhP�č7��)�&��L+��RD��H���,��,[�%t'G�"Bx�j��IDm!�%$@�tԥ3�!�F*�8���0'���`�񔥑2�/��9�#=���ڌ�K��~���@�	�Y�3�d��s���S�Ǜ��Z/D?o��蠼��AU�q}�)G|�h!@���'����D0"n��,�+>`F����3��a��(`����0�dJVY�+�n�	u����-��Y��8A�Rh0w�^_�Զ9']�I��߷U[�|��mh� K5��B��(�W��{orX@Ѥ���M�@=��N�Bq��C�r���2�2��"�A�!�1&�D�3��oGs:�k%����<�1�kr��$��-mL��s�BFl��Cי|/d!`���{D�Q���=��$���T�$�FM�"��ဇ%���Z.Fi����'�U9�E����z�?jz�`/���c���H��ɗ©NB��
�,}�>,�2�K��+���$�Mi��Ҁ�r�ŷ��d.��������:�B͒�|�ڒ�pz�%�3��N��+����֑-aݖ��i�U�lR�P��nt������/h!uF۔�I�Ր<��x�g��t�1���l�[�tr����5T3[;6��F�Nc���W,�!G�q۲n�;�pW^8Gff���W��z�Bڈ��V_�-��gw����Qu'=]�[y�#��ӕ�mЍӀ="�N�;#竛�e���FE��.Gkw�����T����a�l�(��d���c�7AS�˗kq�V�y�#^�W�q�������QYA~~�����a�8e���'���=K*+�e�e�&턪�p�2�j��o�$S.�P�5�_jw�F�4�\���79B��:��L_l?�O9<�-c�_����8�o+�^������0�1��$��6�;e{Օ�}�ʁI�h�AЌ�C]��-U]�&���K#��m}í���@̘��P>�pD�V�z��Y8��8���v
�s��`��ぱ�(�����âQ\�⌛�%��lu��Y��� <��l$�7H Q�����4��磞�R݄M�<߾���	r��e)�t��یPI0r��G~��i.x'YWD�����&'U���&VRk�8�|��b�����V�v>j�I���/(��I8��H%��dt����66�����r��fuLx��^j�Y�e�b(ȇ�-(Ѽ̙��-�Ǒs�W.�C�������Bkb��}�����Ix#B2Vg_n�?��:Z��I��vw#��Y�!E�۲� `Iq�Ȳ���F 3����!�+Ra�㺢�;Ƞ�+�H�ȼ9�B�oƵ<:�\w������.����0�����f��x֌�/�I%���o�U�T�����y4VUuv��6X�8���f��Y�9Q���Y��wm-�Tʼ�q����7gʾ�����5;���CO��㌺�A��="8p��)׀� ��f�hkȼs%����U�P
�_^�c�����/ǆ�1�� OK���aQ2j��;�Ez�2�Xl�urܫ�\T���#�B�AB�=QD����+�Gi/�i�Q�@��z��:W�3�X�ˊ�LN߱G����ᶭ�+��F�Y��u1O����������O�.J@�L��82:\	5mG�_��-z�=��"��?�`͘܋��E\q��.�I�A+�L������LZ�q�_���z�=;>�Q�[|Ns�Y���O�G��Bo��^�+>T�W����k��;��ʛK��h"U����L%\��b�8����8N[�p��i�'��c�,��{.������<}�IQ�:A���}���y柂 ;uD�E<@X���9�}������*�y�չ~$�t��HC ��*�_�8�7$X{��� ���P��l���&�[�	�	����u��hB��C���y��V�����U��]:�z�zXAi���{O�"�υ�^$w�vy�.z�%��N5�P��hi^]�׆�lׄM6����)1�J�v:"�0�z/}�ȑzG�LAO�A�"��F�q��0E�l��n>�[���M}�@�U�y�Q9�ߝ$`���N9�#���)`
����t_��~�N� �̶�/ ߊ���>f�=�H ϗ<F߁��wpp�^��Ʉ$���1z�~qQ�抟K2t�;�뷙����U���(�r���i�aMk?���o,^_WE/٠��,,,P���fZ� �t�<Yq��6�`��n�p�u�ߤ1e���ຯ��)�DG&�G¦���.���d�Kw�9��\59����٣"��:Mѐ�2��b��{�x.��(�A�F�|���Sr���FC���X���T���. UԿ}���)@�s���F�z$q@9� b��ύ��U�r�GM�Q�P����rF�����f�B��k�"�5X߀u�!���Q��_�hҠ���I�޵>F��&���7��j�V������^�4�Z�2КxJ�-��]D�>���`�>\�{M�/&% C�?VSSC����A]�?q(Y��w�~���~�B��M�q�PW���="M7n�[J����0s �!���!ʭ�N
���K�0��^�h9!Ţl �����&-5�N�њ��闿�A��ε׻��m�.pN���~�-o0�(�aRM��ٛ丼E2σ��M.u:�������v� ��OLt��_��]�ew ��� �x'L��1B��Lu˶��ooM+J0��ɛI�z	^�x^��h~X$�P�j��� | ���M����e���-����c�I�=����b���2�sz�vrF�����hVx��avȠ�}���f�l|��A��x����g����o��ѐ���b�8,��&U��`�+V+�i��:ź.��:���3=��n������sq���Q��}j�̞��F>����a��E��ԳH���+�o�p�-K����22H���'�C�I42�H%PH��6.�K�TKډ�5S����Ԡ/H�q��u@���j��J�v����=�rqմ����|Ծl7;�tV�AOO*{�&�Mk�꓎ԯ��>�����/���#���R7��1cS�z��5��v��@��wH4�/��.݁����������6#p�g��k8B��a;�� ��X���r~?o)c�krT?VѪ�Xt�S�I#��������q�����J��7��#Quה��󫽋C�2b�OY
�D��nCO%\���'�����7|�gKØ�`�=���٧�dSO5��</	�$�#����u}g�9փ֠�����s�V ��M'�<e�R��[b��&���,�a���!�@&�U�+��lX2�q���q�/���7;�>�)���v�X.뜵��Srǩ�d�Ū|�7W��[���t��835ݗ�31?�d�{��T���t`���9?�S�� �c�>���{��J�#J]M��&��	��/[~6����� M��Z4��Qf�L��8X͍1pN]e���]���#��ς��#��퓤�h�,�Su�~�������ő�ڸ��T'����Ǫ$|O�7�M�)i*�-))2[�fgȝ�T�C��������X��?
 �\��^�y�W���~���C���W�gb��s�/e����U[#|4ZZqk�/��R�qN�����-}�Y�9���L�(���^�Sp�U@|�sbCO���v>g'�i�YZ�e����KK ����D�����J7a�f����q<�U��Q���>
�D(�-�עMr�Ng�T��v��i:���tZ�i�bZCCC�dπ����������ﺣ8�0����Ⱦth���p��=x������j3�3�{����ܼ�ω	I�3��w�$��ݾ����E�=滽��b�e��ea&�������,oL'��W��*詹KuK|PX���wֵ5}�����MD&�ZD-)��`��>^j3�!Tl�r*�녺��v��[�#��&[[|�p<���$:���w|7�ߓ��$�^�:�Nf �j]��7V�éwĀT5BRvz�G����G��T�󰓚�u[�� �Y|E�J��ӱ�x+y�j�%���8qab��U��GO�5?��%�$�i������y�s��t��Q"/n��^���W5O4����SN0x���M,;~��r)����|x�\�����r�E�͎�����J�rp�s��db~8�.>�LG�7�z��:�ɺr�{�]�6x�Z���swNƫ�{�>�mg�� Q�-(5oC�Ņ�JFqZPɜx'Y�B'XQ(S>�\n`���8g�X0��f�dl#��]z8��i��y�G>((�G_��D����_F��?V��S����1غI�+ӎ#z˅0|ȉ�<��,�8������;b����x�
0�?{MIT��wg�|�����y�ަm����?뎖����?�]a뮤z��s�?p��SuK�r5���x���9!��qE�:F\3����L������k��c�v��620F�+�,ܪ�ό����E�������

*E�׺�[�C@y�X��L9�r��1a���4�ރ<}QD���Pĭ���b��ќ`bwr�6��Lޚv��c�{L�<��}�a ' y�aF�l��B&�ě�'7��K>S'���%��`jǀ4I��2�ّ���Y�s�?��tzo���(�D���{|�>�������]�\��թ�,8���P�w�I`A�G�K��S��a����0(}\�q>��x���8����J,	x�6��5�S칞��}�%]ԫ���#�J�Ɔۜnpd���1�w�Ռ}G��2?{%�������Zu����"�y��`9,�p��.��W�j�?��KC�'=�P"J�f";|f�=��V<�\x11o?+0�㗓4|�p�yj���G%]PK!�1����wN�El=�C7O����}R"N�Y���_�A:[&fܥ�j�E���v�����n��v��5����Q���n|f��^<5�8�غK3��h��;n}R@���7�D/KM���2���XV�q��_�3^��$��X�:_�Wg�d?:_����b�� ��F ��������ב����g�Lx�I!Gp.��0�� v�))�j��os`t}�5�h^���ze�>��j�\P��1�6�c����B&��\���*�(��	����ӿ�5�i&<sf���p#�/����'5
���Զ7� �� Bv�_}/�w�6��`�r����SٸO����?���Jj��~E�gl�6�-��)@.!��㰀��Y�/v7�GV���qҢj�$�D��ܩ�N4�� y�<�:��L-�����y�MNfò�!A�"{��9�}�4B��WT�3�A��}]�c�F���l��D�,�S����i��jхZV�x7�<����vZC�)]:��)��i�gN�����6�3H:�ޱ5c#�	����i!�����ԙ;��-C㒤U�r��v���a���P#"�J�o0��-�b|,�-��m���nq�T#I���\�Y�m�z��5�8t��N$-��
VX�_��L����0J��T޲rę�GB>�W�2h}��w���]J���{���'��rzq�nf��
q���4��q�n/�nN���TZ��߸�p,�_!���PǬ玱����#ȍ@��2�,�и������ɴ� Dk�d�N��a<V���O �[e�!h
��!ଗ`��� M��V|�-�5�����4�*�FjI��/��B��O�o�n"6��5ɮ�B5��<��0|���%C'#c�H�����S��+���0�i O�"	_���̠RG�J�����U����Ȃ#Od~[�8����5ݯrc��я_N?��g?��_mH���Ry�h��"�e���	���!_9���`�[�Գ�׭M��W�u�gQ��K:���C������w��G�ju�NHM3O����ˏ������C�t-�)�6;wh�
=�/�P,��ךdO��kh{�'���̉�X�;9�Qi�Vߕ����v9dh-'E�l����	�.�ۢO�"[�rl�0]m��t4D���/���/)uZ��w��d$�[��s���h\��=�i]�Ƹ�^g[6��*���?��W?0�i�lV����
��%'��W����t,K�/��/�J�S���W�p�]��A�B�(w4Йl27���w�^�i]�o	^�8K���9:x�N���!]��Z�zd��������8̄3TN	��w<��V������a���ѓ���v�
\%�0�$G s���R[��,��S��X��������N+�m�B}6��fs>�s��܏`�?���n|���	e��A�=TC)�:����!�ؙz��&��S+J�~T���뷥�$��Z�<S����NxZ^ ��S����1��Ck��P�fk�y0�S�T��H�\���H���3�6�?�6� ��{����~i���2���Ǜ��}Z�$@Q��Qh����E��#��xf\���Y-4���6���M��
��*;�;}�s�� OF^֜s6�4�/`��q�<��ˁW�a�t�&�i�Pn��L��������퇎Nx�s?Y[n4Z�P�~����:�� ��jf������ϩ�볎�'��8(��}�۳N������RK~iޫ6�E��@SPG�G^�:���A��QS[%�9��d�?�)˛
_�I�.-�3����H�"MJ���O��%�%C
-�C��q����A���ɠ��mPX2��لЇ@0��u�C�NA53��O���S���6��D��v�{��ݰ�(�ԇ��D�e�PD������pE�=������@O��L�wS��)���5�B�U����y���c&���>;
����A�� k����r�7̡�ZH9	��3َ�.�g�ԛ��@�X��n�6��?�+��*FK�@6�˾��y+Z-Ka�5vqΪ��0؈�mw�nyð�=%k#"����H�	��H+z�/���[�II-l�M���	O0C���[-��{�LT/Zee=�<��/�t��V�G��d�����܊YV��-0��BA-u����_kc���h�@��ycM[[ۻ�*Ȕ�צњQ�U�Y�*����[<�8j��J�Xη	M|��ؙ\
�I��?�>�L�a3�� ��#�hf�����v�5�Y����ݑ���$h<�A�|*�e��5=�^�c��M��h'�\�����ն��������DE�i�M����W[��1��k��ze�m�4q�7 ���n�1��Z���^EjD@H�o�0�L��LF�#�C��'�+��Hπd��$: Lp=t��u���ѡ�����0U��z�b��;�#�"F6I�o�W}��傯#�!o>��xG̪��i�� ���ȹ�z���P��GE���D,S81).�m��/��.5�6�'{Ѥqs� ,+�1��X	��N��ԇ/y��\9a@��/�KFFz��ͬR�aO��� o���m�B86XX���J�� ����M���<3g����g6�CV��X�}�-�(�;0l�����[�;uyC�}'��@�LfOe\}���l���Ȏݭ���{XC޽igpT�:��Șؙ�Y��v�͚Ar~��iw;�++�o,�7o�{�]���≇�����I�����i�]���.�_��ִ����Ӂ�@g	��#S��.(��zs�V�v깙�J�C\�@��p壔��h�"���u�$�0���!�����h��@�ƞ\l�����t6檸sg�|J|<m;a� ò���#��YgƄL`�����J�],y�=�h�R�)�;!�$Qj�$0H�[���5}�0Bq��Ͳ��ĊW���am���	����,����y��D��P�����" J%�w�V��d�>*?2;�SN[.��p�n^Ħzf�.ޑ�I����W�uE�r�#n|"̜	�/�p�\LX +�D�{b�v5���� �r���4K���
Q}ۧ�;Xa��D��YX��G��F���=q?����
�M�t��>���[�#���w�Ta�X�,[����ݹ�to~��@��IP��`{�y
{�����2W����`:[�#��JN�~�"v���R�R�N}�Wv�5�KF�p��6��j�V��zl���	����w����:Q~a�����u*.H-�JCX�t��Z���_��R��|�!'(����}J;P<K~���N����g[y���v:_�����4Dx��mZsS
x�H~��=~-�U�4�ʋ�����:}:�P�MU�&�j��8ءc��_s	���1�N-�e����f����k�[Z'쓢����V��� ��{;�?>��%��K����4�^k^_uX�T)&��+͉N %�2<"�%�T�1�L{;���Li��ie��&C���:�U��?�]�������Ry��H?�����Vn/���$q�����$���0=��6ի8������s�Wt�� �sS�_�RZd��=�.5?B#/�S(����4,���SZ�2�}�XT�w����W"�|�w]�y_�d¬gP�]�1�Nc���[J��M�QGE��\؞6/?+�ʢ�R�SҪ���L�!ی���9��i��p��7��{wXJJ2�G��4�d/ml'��'�~A~�n?��:�+9���>֌l�W��|��(���;���~fv2��G�X�K����5�?٧-�{#a�b�.����-,�����,��z;�H#\��n��;@�u�0�ig�b���9�
_߬���D�����t@Ogsxɔ�-U7�cb���@����lրT1>�?�[��	96��>$�3I���W��>�_7�f~�_?���!����D�~����f�1���;��arb�^]�dmO���Ѐz!)�K�Wjcd��ʾ�sEqku����>�݅_������N�j�T�ǫ'7��x�M��L�8����3ݘ��:�����204T˪��,�7a ����.���# +��59��|7ۿ׿7��|8���ؚ���&S�����!�ʅ�0���S��=��I���b�ux.�?��6Y���y����3e��D,�E��Z��@�W�!��`*{�֨k����O����y���7�ki�<�
��"���L~Ú�kC�����ݿ�W�^�ELh7���ý��䚧)�Y����:�鸹���P�J���/���nj.p�0�>�mq�#��.K[�^�ؼ�� -�k���2�d/���+I����2��*��V'w6�_�k���'��B�6���׮*A
�noNhZk-Uǈ�����iK|��]�O$���*���c�ZA\������.=�E��˛�O�Nk�g����5���0xqTe݂�Vyg��tw�N*���6���_6����!�?�x~�!_��ߎ�7�hI��^j*�Y���,����NMS��@��⒒(����2;H0X�ٲ�uVo()o�:}�N�.��Y~�k8,-�SR�ZPoOlM0�^k]ξ�����\�p'9�yu��Okn��o�mR���#�R��Rky�'�����%}�m˹���:�Nw�O�"�l��޲�M#�Ӵ�E:ň�$C�v��	��MS�g��!l�s�������������,���(�ڻ��#v�˽���_�"��~��������Н��W��W��:�U����
�?�����Eޟ��y����(.�\hkʩ%��b�iZ���#.O7��li�'����W���oF}@L�����fr���CE��$�Q}�����1����h�7xI 	��O��z�=�Y}������ё�p�j���1B>N�����|Ōp_ !�k�t*f�x4���)�E����{�%{�p6�ɊDK/�u�=���c�@`w��I�r`w$�p!���N�s�����"�8�eE�����7�# *>5�m�����9���ս��� X�{��C4�a��T��m��!HMMJ�>�W����=J[O����7Pt�5�ȣ��s�����q/��m�����P��L�#�aMt��%y����J7�qfn��v#�䲏�.�ы����K�~���))��]���܁��������̐O�&�$@7��k���`O���yũ.��7g�f�����O���̀Z|�zÇ!'��e�V�Y��4��:P�5:.֭��@N#�1=��iؔ	�:E��#*��lIY��{"�M��m��_�@��jw�A�gXYoM�n��T���(��*t���2�?��⡔u�ɖ���RW�K�'q�7�L�Sd�E�&l�7 5�MvH�ϳSl�\dh	Ȼ�	��z�J$�
O5o,+P,_�b�8(��n)nZt��������{Y�J�L�~�}�@{q\���Ur8��N�A���0p( �L-ޟ�Q> zNƳ\���`~�J�\CQ	�U�!��o�0���0!���3ZwoU]{,0$�Z��Rf
1y��mw�܇{������͔� 5F���-���K�Y��%~[��6�f�I&��y8�*ς���(�\��8S������R�sh���,@a���I��}�C�1 !/O�ZȎ��~��d���J���(�n]A	G˓�%������\C�)�W}Vz硖��|)Ck�R��X��9�1O�V�K���N,kt�U](�Ǎ�l�+��p�Y��G�����.�#IMG&���k]�%�?,���bW�) e����+-��K�ɒMOwjN��(������؆�s;��,�/�ꚬ��9L�t��ф?������x3t�}���{o�;,]��}ź%9��ի{�Q=�HӀ�@�W}��cpm��#ZU�п�9y'���R��� K�n�;b�i�v+6Qt�l�ԇõ$*��}������9jU�T�#�Q֒E�LFd����S�����&̿�|�;�S���_>�����?�)a(û��Y.V���� |b��`U���F�����m�f{1��c��D�Y&�ۜT��j���o����;8f�(��{/�t�rB#���J��y�uo�Y7�n5����?������z?��|{�v����I�vQ�_JX䉎���@�^� q���_��x���"�(�kZ��l��D"�`������
=�H����Y�8q��
��Ɉg)}�?f��x��v���g^:���Wxp��|F"#��B����#4�Bs��b�;�Ɉ�����[9^�O��r>K���i�L_8�*(�Ha�e����;��3o���1�P�����Ѽ+��H�{Y�a$�kOш�0���#r)��'�P>��C8�M3GPd��>�,��X�"�EΨ[�pdA� �p�dJ֨����sG�&�m��~��!�/כ�����ǖ%��3],����;�DS���yg�t���庁�	��88�7�ro�J�/������$+����G>8��O@}o޼	���#�XU��MT��f��3�Ȱ@B�e�[��Rj)Ax,U���WG%�>��N�V a�o��BU�F�q:ӓ"|���������#���C�mY�z�U^AE���o��"�l�u�=�Ђ����]��0*6��=��y�Zu��k���Y�w`�������  G��G�K|���jjo��F�;Q63�����;]��¾�X�0�kePMhi1���ǈ��~�+瘉�J$O�񮁦���;��H��\�b
#�&�&��;p�0��^�Q�����Ѓ��3yܾEs�
\p&�aO���y�E��,]����?|�:d䵖��S<:�;s��t0�'�1��]M������.T���D��i�[:hh�5i���%�,�w����I�tߠ\[՛�����Q�*���g�6m9� ��E9܈+~� �q�7{�b�2s8$���E�{��S� R�>�f2����o���0�n`�ݱ�j��ܷ�v0x�@f-zs���e�#.t{��i	�XM~��)}#�ۺ
�2��I���c��j'R��i�<'|���D�:ߞ�EC
�$�H���Hg+��NU�����ի�u2�K�Ƀ5�3Ǯ�I9��bj��]����	��K��4�l?Z׺�m��8Z���iO푋��G��78A8m����P���h>��W�u��H�a����ş����Wvv%�9߈�
~���]*��o��5f;��(*��G
�0(�>�8󸳺����o���D�DA�E��[�����;�����N��r��A��	q������4YmO[J?zH����`2��h�li��}oIX��P�gG�����:/�FK���@.)��iD�	�2��5Z�Q pM��������9�^��rk�W������j�áV:5��"�A����e��������Ao��Yy&q�d*��ޭK2[M�f��/��nr�@����uK֋vwO����N��'k���ax <*7�^L$�9�<wt���^܁T>q? ϱu�LZ^%�kͽ��YVǂ��H>	H�������o�Iƽi'-��;,�&�ר�p�S~�H�d�1I2//��L���V�l�ׯ�����(�A��&<�	�pS���5�dӘ��YMf�]Wdt�@>�9�E���	 ����Yq:)6b����{PsJ<"���������;^>�a΀�C%������e�����/�TV�
�4�j�	�2�ge~��Ȥ0����[3��z9h��ֿd��J��K~�k�����&$/���
Ulc�z�K���ZR�f×�G�)�m�HdydR���)��t�5�+dsKt@KI�[��gpu�ŝ\|���@HF1Ji�+G���w�lec&�s������TS��Y�0����G>����BL9q�F�.
������ܘ�8겮5�z������:~��9��x
����z�j}����>5��ܟ �d�������ֲ�ݡ����T�>���7��D���r���߬|q��TvI�����U�h�n&֔&���S���_h��~X�p6��ڵ3��;]���şT�B�W�M��qX#D¼ڎ	�*�2�N��7����,X`��vV���D}� <����t4S�Vq�������w�`��í)p�A{��:`v;���.P٘���Յ�ܩC�4�5Rh7s����3��K�&/*T������+dqb
����4�͘�#��U��g���6ҷA�x ��"ex�M�!//��rO*��(ض�}�7H�/{Ya㨯�\Y��d����剋rF�f,���ڊ�⬻��Mo�֮�`�=Z����1ZKMK����d9fk�'�{��t���z���/lxQ�@A�i�$����n:���R@@rh����\����~�˵�;s�=g����<��;w�[�\�����Q��͊�{��f��vP���Nk3���_h5��A�#x��~0��}��S:���-ϭ�}:>u��	I��ZY\�K�T9N�3]=��`1,E�KR^�$"�[�MSI�>�=�����ˊq+�0����Ϝ���F��;	iVVY�6���a(�3*��̗��W���$���V�޼(��������]\\<�l�V)xS$1|�Au�e\��ډ/�)�<��Pf)�^3��#c����2i=���x����h���5����o������U9��C��rí٧<	ݚ=d5؋���qNB�qI;1�M��������C5�٫���ë|f�ǹ��沑]�%�YYXXX����l�#�%�s�����c|�����z�.hF�	\�
D��o���y�f���:-���a��4�t7�:�y���;��_�f��K�[]||��' )���SͳY�M��$��X��L?��� n?�9��0!oY����dG���7)p���u{nRz:�[���s�������7R�y%/#�i��!�Sq6`�����CZ~c�5NV��:
�0���e�cP]0���i��w7�;BOv\:�_�����)ww���S�2�m�p�l�Я,�룦��h�� }ۛ0p�$ŋ�;�[��x|k, ��r�Y�D��3�` �f��.�:USQ��`\fcnn�IuF��8�鿆�5�x�`�
h�1id��>9"�^lzt�=Nܽo�Y&�����:qC^��b�GU��3�K+yyyy��p_�y8�����o!���<)I�#�M���mcK�}Ĉ1I�C�JMH��`ܒ�#��3?g�,++������߀�_�z@$[�]OyD���j�l
�X�U:湩����gs���8�)�`�e"�υ����iT���a9w�� ?I�0eפY�6��v�j�?����'��_��wҌ�v��!1W�88�,���������=t��@~��	_�U5�D�V�3���M0�]�2,�_x\��Gٖ��_.u���r�]�ttt�To;:�N~�l�(�PZ,���P2i:����X��1_��}���ei��^Yܾ��ƣ~K�fk�����&�/9oK�!��~�f�;~[Z�vk�E�*9K�\�؇�iksJ����T��R������=�X.��
��56��n��p�-EZff��MN2��_��O���o7YkD�t&�^w�����dK��G�s��&=33��3�%iF�$'e���@ͼ��#��x��2�E�MP����Qjڗ�S6L�6�Ћ��$-+;H���� _�D,���ݤCk>U�)������<�tG�FG�	]�G%)�ȧ��U鴞gS�1�$�f"uyQ���k)�OZ����8d�˶���D���2mG���v��J�Y���v���<\��C�4K݃^�S�º���f�2����V �%�ss�6Ze��+X a����?|)�I��N������z+be�Ne���;�H/�r�LC#Y�~���ԭ���r���]�"A	I�>�q:�:9���6��_��+sk�K`���l�':9�����~������4&� ��7P&��/���5$�An2�ҙ�{��{$H66��N�J��Ju��%���
�F��:�VP���,Cl@$@�_�;t�r�t�ф�"�����q�Ւ<<<��K�6������M'�?�)�����y*��͊��t��o��)��b�T!2�92�i,�B�|�8�f�������Ek3�8�c7϶�:���;C)-!d�Мd�C�M+2]�|E=��P����~��}�`3vJ��27Ɉ��J>ַ��L�N��TH�,{��"��R�Խ�kM�Ɵ�l��]�ډ9y���ʹ�
nA�?��l7"&F#s.0(��z�[��v�vs�Bp��ݬ�XO8�~x?�|6P�,����\�>IM;�t¿-+�ʐtX����@5�5zx����*�F��7�Z�� ͘O�m/�_�W;o@���zߘ�p���{$�'(Ԟ��fg?r2l� �*�}�ڹXZ��
��3,YYI)�N9�H���P�<��*d�N*��9���'R�;rCHy��
,�p6d讉�?�x��#/{w&���ﬃ��sϋ*�nW��f��5.���}f�֝,�|�4�޾�<l���_� �l.�m/>�+ӽx2j�QZ l�;e툗�v<�᧽������#ъ�T)�v+��]�hF#
ӈ��r��~�|�uM����d3��º�v�Sj' ���O�`���,�m��a9��57��6�v!�X�;V��+�"���jS�F��t=�;+F�m�d��U��N�x�x�>��$"��JG�i��q�hD��+�w�>'>~��R�t��sʳ^%F���(P�-+�	n��xU�� ���έ�=��%��� O@kEz1b��U����&]^w�D=dz�p�� �FH��wœax} ?�bp�k���U+P0`�w1��eF�Q���.�$�ߪˋ��IZ��������YY��^7��R7���U���y�~�!��_	\�s[2*���зƈN����JJ�GC��mh C{��U��/�eo,��v/� N���V�R�:�M��H�p�1L�f�� ���DJ~��Z�+I3�����T5t<�3��?���Qu@������,���;��s�0�TSf;�L��&*�^���n��	&i"�j���͓��%v���/�N����� ��>Ɓ�>���;߮�Q-8��n�Xp����_�Ň�nl�齃ͩ½�=��(�n��J�+I����{��u�R/FӢt��pi��'8-��N�S�|�//N�ʌ�ت��^����
���du��ǆ�SW��iT�o�Z^����I0%j��I�I��h��n�:�{�ѳCH�$z������\��g�~݂L-{y�1��6����z߯#w�hhЧ"VIu����7V�nk��=���.�~���](��dG�!��%}fu-Hi��8�}��Ҳ�Y�t��}7_�B�6��j�D���߹ž�l#�b<���>���Ow�/�h���e��:��r�%��Rv���"
�Py�7�����TÑ���y4p^���O?d�q�;`��#�:] 1!�_�������E�А�8�+b�����.7ż��x��m��q_��ZҊz=*�&�Mجpwn��PE�%{bCs8.��+�\��}`+���x҅������9��.@�I��~�dwa��</�[Wtb9f�))��r�L]\׳ж9�D�!J/Y,3��{��W�=چ1�h�H#�v�Y�H��ّf�L�r=G�.�ucg�~
�}m�\�%ewr���#�c[�$��A�*7������i}�͔
�CL��&�e]��� s��w��MV1z.��k�E`Pg���|�M�A؇�����(�Ҟ��xK�����*s��Rc�>�D���ն� `۟�d�E>��:ֱk'�6�m [�vؘ�H*�'-����[������r=��2$S]�{3��!w	�*l
TP�
���ǀ�|��ݕ��㖝]���G%d�Ѓ
�%�϶X.��6��L�/��ͣ��!���0A��ђL�Í��4��x
�vzz:f%�p(��"<&��_����$�v�ׂA�L�o�I~�a(�����b�/�*�F:2:�*�Q�����1&�p~,�i'&R�����XhW��[�W�0b�Le�)ϊr�����\+	Γ�aA��=�l(��te�z���ߤ	P;~�7I%���6-؛u����Е�$��_A����8�Yܲ���^���!D�$3���y�$����HmS�X�� ��_���	��I#�օv�Ӭx�??�%��[�յ�Ԋ0�?�`�>�>��R;���V�����Q K��Հ��'	�Ɉߊdh5�b���nzY0��X���"q���ޜ1ݙo�X�L����S�^��&����Z(;XR�M&K�4\Zi��8@f[Vj��B�=~�@���p}+f~i)�)��;��3�ks�g\��M��H|
�?�EEE�
]���<d�\����I�>\J�	��퇌��o7���������T��7���q+�5*C�q��` �<�m�O��i�J��RO�זǂ|9 �?>��:&�NI/�Ҳh"{��T�ȶ�`ӕ�z��A�mڶMXn;����B�׮�y(B?��8.:g�	������ΓWonݺ�aH��>�5�*캈��:ۋ���%�ҍ�IV���� 
�����6��I�ĲK���]�9CxlS{w˩�۵N&M(y?o��,�4�_�e��9>RI����dP���a*{��?�����j�^�SLJ҄�쯀�222_��BLp�j�m5�d��;ۢ�J̺B��y��g]��G��נ�v��T����D������3,l�@K(#�YoZ�ؚ�/� �2 |�鐐0ʠ�Wxnm<%@��"��2����??a�O3K����/D��s�L��Ɉg�8<Y瞫^�k_Ei�@c�@��m�4_�N��`���� zU.H ]��9�/<��((4�%�ɞ*�sD���XSH����f#L��j�s~��R��M�ᛃf5+�&�V�hhi�BTi���,��IE�8��6E�ʈb/,,ľr-�c#K;���~AFE��p�*����G�벯HTWۅ�l�K���.�]��E�e=���X0���ux��:�4���ϱ�q5�m2
0V2m؏�;�+,�9��[��##�,&��$��`�.�x��[��q���[��e���A�7\����e7CN�A���.�5������j��y���ͳOr��ϭ�D��feI�8'8��(�v��������$๾���
�X@:=9m�r�n\}Z/y�@	֘M��u���a�!������S\���ذS���44���&�C`8***����̮�J��r�2F��fj�T	�.">>/�J�cua�i��8��V�����/��]	n�^�?��:���2�A�^�����|�k%l.[Ӛ�7�7�ɽ� � ���0������Oy�Ýڧ>�O$+�����x�/�Sb��;�3�{�k�����ґ�f*X��}:�;�ע7IHJVV��i}��J������W`4
�&4"p&.$PlvX/t���5J�)���]٘�-���>qrLj(�����X����֏������T"xd���.��_����m.���>>��r�F,\˃إ����!��h�Y9��a3�̅@:��>���2�V5⧊�����D|1�_W�u�/�^��_.:�\��b���L�Ut���Pp3׬��%�@|�������A�c�� v�yݩs��?O ����������;}��X,�����~����gmA/��<���5eҫ��l��]�>��a``�D|����#6cS �O�l���� ggg���%�NVr���+���;::��5d��1���S!�	[?HL$q�ǊW�6e�b:��NL�f�U��C���d{�캸�ا��M�]	��~JV���l�D �D�[�َ4������ԠUT���'�����o$�[�4���@2%���Ӈ��H�> Ł�D�� �aY�]s��>p;���Sk�4r!��&l��^�j��u�4��s��q���Vc��Z�}b��;
M�w��3 ��r�@qu\f>���ʊ�
t�]��t����MFEFf �[���Ga��a \tٌ���f���A�^d�����Ɋb�QΔˠ^�ޜ� (H�k���҃f
�Ԕ	#�U��rТl�pU_�.ce� vv���%��6+�*�ܭ�t=�?���{Gu�;t����uL��<�wj��M��!O�R���y�.)��H{\w�/�	wZUڜ�#4����(4yq�S秢�S9s��U��R��������r3�b�9�^�V(E��.[o����l��9�����L��\kv�WV���Ӽ]qC�.@�I�؈��]�%2�����I�9���FO	���4�$�ؐ�b)��!+}Ε�����L��'���1��<B���>zm����Ҹ��ې�pk �I<-�B2*������pU���n��Z]��S���7X�l�0�Ӆȃ���}�p���,1~��&ۖ�b��]��V_�y6��Gi���{A�,���I���*jj�{�9�WA�^�wKU���0�*D��ӛ�X�V���d:���>K�e2�9^�ڮ���LK�F�����L[\4,V6�Ӭ�ˣ��.�t����y��JJJЛM�N�:��D-c2�4�?�t���|�D4�	�g6�M��W�H��QV�~L���HyY�3�e��>��岝�P��FQ�Go��xE����8�}��>�1�9�}yN"����Tt�hI��.���j�s΄*.�����	zl���_,�o��=�;�6�sP��V�]������R3�ܪ�01��d�h�sE�^o%/1���p6e�{��^���Z� �޽��!�R	�?`e�?c��h?Q�}��XQ����L�C�?Q+=x�(>�����glθ`�R��{�{�*��4����PQ�ZZ� �c+�Uj8[`�?�}���7�יK�v���x�)ԇl��u� 3Z��:��ٔ��ٯ_�F� F[W�<��1�߈)`�X�� �;i��6ڕ�5��q6�x�z�蟿�*��;�р, ���.��Fݡ����0
�=��N���#8���Oxd9<�Y6S�s�'��������Oe�ɮ>⫿���שiC|[R���*�{�j�/��/���� �`��Y�dŤm�w�E�c��v����ѫ}�c���F�	E�q�I	$@��N2�b�%9\���|{_�B��tD08�|��g����������u?%L�>נ��D��^�:�1R��fs{��Wҭ�ԝ ��m�'�5���HL��R����o���BK��������#Uճ�BH�M��|���8�z��w�cw�U���O��:���-��UX)Û�I/kBBN6�k`0�:���T��}�(���n+f��kеi8/B\�-��f���*E6)r숖�_�Y�2���e6�]N�ˊ�;ܿ����'H�9����L~�zv�0^�U\'��A���B���#�ٰ�f�[(�S{T��J��/M`pp�Ͼ�� r�����w/�H0CJ�s�_O�8Jڤ*F��3\�Ny&֯���
M0|-�n5�ԇ2�}�Le��q��x\��O���2ýe%A�n�g�%� ΀��M{)h�����*:�������pA�hY:�g����p���(������z�,f��E㮍ZE$FY�o(Z�W3�_���) �g�͹��bv�_�Pt(-<?Ġ2WA"�T(p������6JEc�j.3��������q.�5r~��g���BpV$[vU#�LO����cv�?��䀓�upMy(���\m�}��O���Kz���9������&�%I貳�o���^��y�_��{����ޗ����P���I�SM�R��7;;�� ��i6[�F��V�:%�xTE_��[� ׋7%+���������}$Z��,:d�ͫf&�X�a(��#51(�v������;�ա��������6hyX�}�y�TD�����i�j>z�|~\��f_�����Ps�㵴�ą�p�+�wu�� di���k"	hMU=��m+ �z�O-����<OO�@+7�6ai�mf��T������F�+��ۦ%gA�;��Q����5"�[lt#۴���ds���L�-�B��'\ NY�CL��Gҹ�SQ�-(d���&��ݾ�iIfk��9$� �V@<�Io��*�$��$��C�%gW�J�.��dmtP��	�	E^Rߛ'���H�$2%�=��r��hA����4φһ�r-��߂�P���l/L����@����0Dn����y����ߨu��/'ŸC۲�/���9lG���̻�y�Wrreڸ��	"b� �8P^BM[�X�8���bͯyN���[N�w�;���]j`
&_lZ�{z�!�6#�J�Ye��%fAF!I��9(��������H1�׹�Փ�x9���ק��Q��4���y1P�,���8��EQ�6��vu����ֈ���=��qv�x<�q��ԢFSa��ֆG��2�DvG�3�^iF�0=����we=�{�?�X=��}�>�rhA������~\lV-=126&Y%�&R�c��	ۻ�biӫ�>��i�\C��5���Ӟn���P�6X�o0&�a�^���f�\v��� C�YX�jߍo��|a��nT�d�$�L?�|��!�f�h�çRʪ��		�>\]?����likε�D=�ڝ����!�)�xթ�~0����d�V��8�b��P�/�QQܔ��Q� Y*����Yl�3���h��s�,Vdz'�']���G�5K����]�K�9��s�F�*@o0s�C4Q��m��|;��h�i�k����S5�\�p��mv?n��bG8]�a���1�)�G{�4V�|`�ܔ<�JL^)���䴊bVҵ����{���~>ʚ�
&��-��$˃?�ǅz�vv�	�<�G����dXM�OƆ��>7��nA>�vS�B¥��2�K;�)�!ߕ�%a��4�<�K��R�s�g^&@�S��	^��S+�w\�����"���S�����w��V��ihd�����ܴEd�O�\{
��>�u�����/M��l�����ѽ #�$�����ER�`&���b���$���{�y�릗0�O�ޗ��ـ�Vc2ℇ2�W�����*>���`�^^�}<cw���B�/�����[�f���oc�Tg�G$?r�m؟�2iV��Q�=
��a�e��6!`� ��Ν�Z��x+(q��C��&߯{X0A��N���˓�C��J��l"?q��WӨ�u��e��F�:y�0�z�-Ŗ>Y�z�����WC�����cFA��/��)W{� �9��19����6PKT#<�xf�Sw��9�q��0w�;V	�6	a�]�D�(f���ϱ��9��}�����!ߡ�0X�r ��^��t���~����f�`r] Yɰ������FK{��%�I=̞�}c�v;1�l��rq{j�|?6pg�e�Nd:ք�Ũ6��`�ﴴ���:�yjh<�K�Ca�ښ��P%?DǱ`I?�A�d�?2��e��Z=/���)�a��	�����[�B(E��m�ҒӕF���)�]���{S�hN�ȍZe��_�{-����_�3M�Y�I��W�_n���Lsvvvrx� ���u������H
���E=v ����>jy"�$/����f� S��!o��@�zXVi� �ݤ̷��#�j `!(�d���R�B�����3����ꅘ�w>���Ӎ�</IBW��~��ɲH�0`���W���QҗG��Ř��v�����N��Dbk�ð�蚼߈���Z���Gl�YΛ�+�%�O��X!RCH8x���eLTڙ��ˬ�1Ϭ���>d������s�s�9I�d���S�~}�8�"GY����f?[�D������o��ي�b��H��_X�L�or�����':�}p �Ğ\*������)��͆K]��JF�ccs8�ƞ31Ɋ���m�}�FSgg�j�އh�쓫��c���J�%�J� 	׼�Հ��
U����6��F�ʥZ�����6ш�?^|l��]Vm������2	o}��I��]����L��?��a1���ߋ�����/�`	�1�=�񢏓uE�F�U$
Cz1b�%�q�����}��w0��g�J�Ư�D*�*l[��f����bc@'@_�x�cC�$�=�B�[������{a5��5�o�l��
�ue�#u����?�nH�DVK�8���(!�D$�$u%��;�U��������տׇJ	�o����Y�oP>�$�%�fۮ�,l�x�y���h�ދ�Ah�_�k��Ž�j�r��6T��x��Z`rN ��!�������R�>;�L�|y0!������PT1�e�ff򣇽o����]�2�����9��u9�Vo�omZ̝K�(I��+�
��'��Ԏ����e]O�*� �O��qS�/�`���W;ǯ2a�Dw���쒁�'=�c'�Lc�f���v�eΫ�j(ĚȠ�wx<l31�^�n����
��Q?ؗ��؞ڤ�_\��RyĎk̽�P���k�PQlz�b5/��<�3��w5�CY,h��Tu��/�h3K9�a���|Kml�d1���㛥�exk�p<��I�P��>�>1��I���0U��ʈ#۔�;wb�SEhQ|�xۍa~_��.���[<g��U��G^�O�X�P�t,����}F�7��{��-7w�7��Hʴ�_��D�f�?�M��fP��f��k�J#��;����T��ʴa�D2ie��e�ý]t�����}L���)(ã�eı�
���n-,<�B��Q>�v�������������0��gX�������٠����]�n�g��O��aw��L�|��?�j�����e���q�����I�h�I������@;B&m��i�ҒQKh�Z�o����=��QB��AHHH�Ĵ��]�.�����@-�9n6U_�Q9���KZq�p��L�
��e>Ĩk�ɥ���n>�.���dV�:ݪN�7*~�;��opn�_��C��59�?t����<�Aw�j�**];9܄�J�C������&���ʛ$����!,
�Ӯ7�vu1��k��w��9�ΐ�B��H�lmq��|ǩ���,CU���h�B�S���x���aLNc��������m%X��5��Ru���s����n�<���2_�$�����k�����NF��)��G,�)h��ݻ��D
¨ġ������Y�u���=�Kr�W���'J�{�L����d�L�)����9��y{��nW�ͺ���(�NsG�t��efb�B\��x�<m��_���L�1BZ��cF�=7�s�7������آL/�O$��qye�ٰa��c�f�Y����س4xhAԾs�D�loo��ׅ�E ��,	�� 3ɘ�7r2"��i df�'�B?�7���Ru�ߓi�v�FD�ǅ��< z2��9�:ƈR�X�ʭ�Aܹ�7�$+�}�%Vy�4|��p�24z^M�9m�㸻/�T��b(Ӿ��Q�3q��������E��Ri�x�}�ܶ*O#��Щ�U� ��ɩ{L�C�"�#��@q�Y���לϧe��֧O�&v`��z��G��/	��(l���f��JeJ�
_�Q=�P<��
���|�e�G�62,��m��6��>`|�h~I}���2�7I��1V2�aԸ���{Kꋃ��A+����$�|�t/5��.h�J��ю�������P%I��b��w�:�����I��n�	�:h7ɄP�Vd���9y��t��L[.����p�\�ˋ����B�c~�C�����,��� ��D��s���J��wH���l�C���]���T���:���+L�{F �)~7�ͻb9ƪ21��?����V�0�o�C�����
�5;��6k�a�����@�����IC��bˡ��,'�M���C�cՎ��7�F��7�;�p0����,+.�7���ڛ����MT�Z����9<�L��z_�(HXĥ�<�-X�x�Ο��	��vh�yS�
��gT�&�G��m�����j���e��!� �=n��/Ie�ZfD�����,-�� ��n�ً�;>Y��7����%�Y[r�YW]�Ǟ�q�*�p��� `�;)Y���`!:��?~���S,#��<O�`�ܵS�;p'�oy���/�O��B�R��T
�x����G�"�Y+�AÑ�gI,��Ѱ	a�v&hQ�$��Y�I�,�o��~�~��,��/�,�>Y�t9�o���	��@P����R����q����;=���2�4�Y�9J�'�\LP�Od1�_�L�6p��~Ϛ,I�<�^j9O�����O�AD7oE����h�	:��	!��L�x������"��?�F�BFG�O�1�#3�W&��>��@��֗���
���������J�P͈I�qc�����@e8�+�28�K�>�����@�SD���>0�>v�	!x`�������k¨Χ�Tp�1mf�x<���,1�Z��r06+d)я꺅=�/IYY[s��׭�!�8Nl�����сJ:����d0�,������k�)IIj�[����;?�NR��2/�݌R204T��,�:��T����vv汰��@K+շ���w<��_���Ʀ<::j�K�2/a���AF5BJ�N��7��<	r����ʙr��:!��H$2��W
I)		�/i�VY���v��v�=�,X�V�۞��зwp�SKJ~^IE	�{���+'�{Bu��	�`t_#�����D���x�T<1���y�&�ƛ��o��e���~�����[��	ϓ=E��@���\Y�7��#V�K�u00��-?�!�ǜYE_�L�mL�u+�����Ϳ�}g3^��y�L����_�{�綗�3��w���שQ����?YaXG�J��0�+�#��9�r�ue<�Y|������mJw��)2--�0#y0d^���;�ce[}�C�3�E�˫>9�&}���:Ĳ"K���p�K�R]�5Z�?�����P��:����i&�r5O�W�jj
�9Dv
8b �8��!Bՙ.�w�{����K�� �_��f�� =--:DՄ3NV��Ŭ��T�F$紞p��(~�~o}���V�ݘu�*͒�����{��]���pH�~Ql!�ǉ���I+�]����Nh֞g�|�k��2�ًؽ�����k[��
���}!N\f)��SߪcXd؆=Q���3�"4�T#+���I���S�t�W	ii��Nfna���Ow�:^��s���2����v�v.s?�F��t�9QI��d^��ϻ��m
�[�I���a=�:�`�t~ϓ����N��\w8���qPQPx��#���G������z�����q5z��Muڑ��2u���G~�D��^�s�FK@<s���9d�E��D���0l[��ؚ{=�ሼb<?T��Ԅq�w�m�3�N&~
��*�?1G{��W/��ۊ�?I��=.E`�����æ��fW���w[l�e~��.�G���������/�t�TL��Z׬s�o��AU45s O_T�n��>���=:y�Z���I@���Z�d��PMp��ӻ<Q��(i׳ϻV�"d�L�\o��O�F@jwx��md�ˑZ֊ߞ�ʴ��HFy_��ϑ_�mR-y^��g�q�8���s4���i��V�-6r�8^ڿ8���l����"�>���*�{�����~�wnV4�_��
���W�}�ͺCz**`�,5E�d04h{�o!D�ٗ��i0�0ZNN���п����O_��f}u�*�U
UTX���]�C�'��7��y���_zF���|;�(]�mQp��};p(�s������b�9�b;��.V�IE W�5�̘S	���`�9�]�RE9�<r�<ԝŌ�**YYYJ��Q���¾�b����)��,3"..��5IT-`��;��w
[�UA����V��t..'k:�ƿ�\�!N�2��liy�/]��7sf���v�z���d��u�ޒ��ГsUڙ�i��t���#�9� 89���!bG���EF;&ڂ팳��
�ll�����.V2��h��v+����Qx��x�s7�e�33ɽ��@+_ �2��Ó�WC����f�b9�4n�噄�To.�%ɿ�,�[�t(u]Յ8?8��V9��/r5�1ULPf���;7�5e^�nV��ic�����DN@���ARO���Qb��Rw��J��s��]�Z���ȯ_��7���Ί�R�a#Y�
���X+�l��|ì�W�û�A�GM7�q ǡ�ݶ����Z��I��,���R��k��V�l�����)Ӎ��A��2����7�.��b��f����K�y�լ�O�@#����df��,������Ow���v���ӧ���蜩ˋC�Bra�Xx�;<u����ʛ���� ����888ޝ�ݩ�O���׭&k5"�>�]
^���Cί� w�ј� �B����{�u��EM��![��x� T(=�W�sL�{�����I�~�<��4n����_��3���ݍ�1�HH�Z�ڎ��b�?�����H�����k'Gs���L��A���>��&	��NF��rX�{_xt�q�Oy��z8b�J�&�:�*�O�}I��e3t�U��˞�����|����������1�7�^8P���_hp ����3d�յ��z�Oev�P�X���|m�I��/�O:����n�("b�<Dg��qb������I�,n'�L�F��uuD�B3���;��~cz��c��P�Y-lЅ��fgg}Ǧ&��{_��"�N�DMK��޽5KvuK��T� ��]���~�ܛ����hS�;�:�X�����;x�Q����0x�0pN?M�� �����n9�C�W?��.�\�2���M�Ú$&��M\�����b�L�F��+��}��ئV�0)��]�m%;Z�Pu==T	��]z�����.�o9��K]_1��o΁YL�V]�e
�5�%�p���hJ�����-AD����������񚯍� ��V`qzgb��Q�9��Q�;$��{+%���[h>��^�L��W����⠢�!U,T>;�RـN�L<oz�nX����2Oz���Ǎ���Q��"���P�l�+S���w�E��}����'�N�'�C�Ӆ0V×=�����i���K��Q�s���+��U�eݓ�O6N'�,��O3��g���8��]�޼~�� 6����GI�σ���|���E��MEDD(XX
��L%����h2��?����-�yttt4�ʔǝm�z}o��d�C@i){$�N �â���vV}��3 ��lみ)�0�%H����(�!�}k��ߥ?e`���<��^,UH36'AWW7`lLs`` �2�����9���$�m��|�*W�ߧjbc?m��f�XR�μ���n
#�����WT�Q�����FxM����-^����	����r펎�&\��y��c���|����Ç�999_���C�(��� Vɒ={/hz#+''E�Ʃ���h�uFQ�^����9}`PP����8��A���P~99���$9�� ����!<Ύ�C�S)��ji=�ܯ����3**����|�ʁvvn��F"ٝO�*��r�h\�K��S[q�]<��ǰ		�6�c��Fs�IZh��щ+�=
��PTQ	������Tt=�oV^N���{���?&&��|ii�p��u���9h]c��C�g�{�o|/nP��b``�{���ׯ���؃���wXK�T��Y�V���T��酳#H��>]fjku�x	����MC�(�a��o����Ⱦ�i����y��H�M]]�Λ��9S���x��7n:����5 �#��8Q�,����ZBJ� �lQI�_D�\�U43s+��ř�_�(���6��|}�ZXt�x�rB�����A��u���YlԹOEG�fҽU�&)y���AQ[��n�/Oih�nݺ��5�^.���	3331��ۺ��h�g��߷[� �� >ܜZ�����I��W=��� vB�U�LQ�����Vj��˛~�������Q,�}�=���ʃ��7�o�� �5<'S� ���Z��O����vTF"���ǿp�3}�捠�n}� f]���t�<l�>�E�/Ĭ�-�-8��q,�l�ӂ����[�V�,��e�<p8|��?����.��)X�Ò11q��ίqq���m -,g�RQWW��u�Y�O4� ��Y�����*�����-!�YF_Z����Պ�0+繠P�~�g����PT�9���(<��KO�Q�����'�kÅ�=��w�İuv�:"��͔��=�^H4����u��g���Ӝ����u��U��r\}}���<�Ճ)(��$�8��hVл�_�Qw�鎹E����R�4�T&���w�t�󷂺�a!��kגӨk�UUU��{���D��t�1������V��=�V�⫎���#$��{xxz�ln�����{ ���������'�뵵�o,e���tZ'�c=����S�2S.����u�ûw�>x]]:?=i� �W�	��C��7o�������>٣���Ĥg������K2Q�_��:�����w9��������w� ����-�L^�t�v����M�W�H������ HN���0pvrj���[]A�I#����}���ё�`s*tz�������*^�5��
� +�丽θ{�~��`A���BW^�rű���S���e�:`��Å�
W}�z�'K���z�;#�^���-|�@�}%����Ǐ�<w�98C�"����݇a/Rr��D\:(���|	���EvNN��c��%]����H�=~S@�[�FKf���~^[���y��)��0��T�D%W����}}������?T[�()�g��,����ަc��(�Z�3r#^*� ��|de�� )-��<�<X�{��ؒ;���8�Qo'W�V�n�>gd����xu��?1��!��|�[��~M���Y��%*��f�5�WO-���y��#^�]�?{���� ;�����{L���m��K�w ����
��Km$d
J �i9�C#��1'�����{:�3V��'''o����;��b�`ep��Ur�~u�`��c&�x��y�<O��ǵ�Xvk)�=�tq~�
4ԛZֳ�s;L��܂VGv����p���C��WC@e����A�Y�͇@�����h=������En�5�r�N�;�nmm���R���y_z�{��f
n�8�}��'9yKN>33���'ܑ�7���?�*��^yF6�� �G\1�)���B�ů��IX��1�!;C,�V\�uz7�9?�ʹ�����+�h�[w:�������ldd|���^���������S��ן��TPT�� �����!E����$��P���W栵�j��.c��D�7��W��
p���x���Ӈz%;�Z ԁ�)))�:,����5�j�m~����{WA(�'/�{���޲yJ(�|�m�5�����9kݻ�)/��UD���a�-��ڢ�oDDR�Si�;�F@���[ZR��[�nA���.����~w��1�@9�{�5�|~�Zs�WNܓw���M�W��!ו��9��0{{{_ʽ)c��_�rs�"����]0v�������`��������U|�"�����2&H�0 c>�--⊊h���bq+I����o�5��^ ��qDTl3��=<c��U��`�uу�Q�f*t�����������9222�P�A_������z!��o�q���IHPA=�v�N1x)�]�
�VSorT%��	��W����,j���W��2�1�})ﺚ�no��#>� n?@WIS3z����G1������	
���X�L�𴴴9�̍--y��G�o�P�:����-���cF�z�oN���caa͒��V@����1�&V�9��sq���Ē�[`K}��w^�UdK�����O�/�d����fF�xz$"���re{��d���Z�����`��\I	#xMMj�ގ���c�@�����Z?I���>cccb�ݚ�"Y��7��֌=l��9�:��Ѝ�/??QY?0��*�J�~4�54�+�Č�i�MLBbhc#wjhl���?�����<��@<D��w�g�(2���jpCCCbjj�NNN ��׻e\��=ܭ��YW������}�^%_���IX��*�^�G@�~��0�IDD��MM��}!��3��zH-���w4��$�;i��m��/ ׯ����).�R�}�0,:������tP��7�@���-B��ha��H����^��2q-��"]]]%%%@x���]]N��xx=�����_ss)�����1�R����D\ZZH@��޼������upv���ఙ�z688ݤbZ���E��Х�bb��}�߾�8r<j�F�IO'!�
.1熁�IRC_�B���rb:u���쳞`TNE)]��"���n~s���H~���`-������=5-�1`{�;.�y�x�� ���333A�L�|D�}/+㊉z����勠�� ,���A��t^,���Յ��F�f�鰂D>���*����C�p�'x�U�P��_����h�hI'Q8�U�� ��\6�����>`��98���B�$���i49Q����g���Ӯ�Y�	��W	��QP6�b�8���3�ccŀ�]��E��ëǡ�_
�\Zz��A>$%� ���3�7��Q�҆1B���~�pk�X|�@G�B� (&�Vd�߿�LO�֚�� =&tv� :8�h`�!��%����,�LV��r������z�" ��==MWy��_��+�P�]\tX�|s..&F�)mjj��f�v�4�z��v(�*'��^^|�y3�(	����Q������iC�����������2�����F��8\888r&�h{2�?�;�#�j�9�x�^�d�
�ߒ6QS������� �֞��(�M���%�Q�L@,9:	����O�v���Z6�?Tsq�&-�^Q�;a_q�V=���L�U�����!Y'yw�FQ�ฝp�����	����x"RO:*t��Z�[���+PTrVjԚ�*�����A��Ĭ�9�3�͠V���r��I:]�M[�U���JU����.v{��L;?=Ө��\��! �L��h� ����̠�����Wğ��(iW�t::ɂ�su�7��o�k:�χ�fCQ�f�PN"  ��&�3jq��U�4���"�@@C3���3[M�.DEM�x��$S#���ݤ�e�b�o��%%]�Jy�]�����Q� c�����R��9�0�����߸��K
	yqppp�PO�0�5)-^�W@��^.U����k`g�Y��J�i���l�5�'�B�*HWF�vy_ )����@�>([���:�+#�D�P���x�{C��wv,ک/\�Vw͂6�u�M�y5���v}-�OdI������G��(p ����脄��ZFff 8��"ܣ#�e�hT<��;Z����\	�󏙎�SP����X�$$$��&����Ɣ���}yￌ)����J�w���Ώ�/��C��Y5Ȇ���*�@ImlnV�� (窖ƍ�(��60.����,�9.����3Y�:���ݏș�c���scEV^��!***��EE��"�AD���m����쌫-&�VS��l���$�CIl0un=�Dv��#no�@��R��R�5�<]�����OJ2�=�ܙ��w��1z�C?��N��U��X����Hdf��X%��<]�2ݣg��D�Hd@1щ��~g��]��@��^�x�x��P�v7:�;\�|'��3ɋ��6!��R	.|tO.���߉�>Q[9�+®p�#���[�:>�bcCO���q ߴ���iu�D��"`l�L�#� =0�X4r�M�0���U�oA����0ͬ�O��诘u��G3�������ׯ
d���>�����P�:�mHg*���"ꈶ�E#cczL|h~��y�ɗ��0���?	���� )-��Ԅ������)�g��#U W��nۜuutV��1���־�����:���n���>�����{S++$�r�1rc@%��<7 � ����먼55~U�^(gW4F�?��֌���w!���Xá�[�P��z�
�$2򋈁�1���eZe7&(��1j��J��Y! �����st����{c]��������w,T�;�]�k�p ���O�=:|�qQ��@H��]@����Q"7X���D���'m�###��q�io�M}����WQ��#I���CW]g9�
�J�95u�-��� ����<:F@'�A�������J���M���\�)��Pu�[����_H�S��h��:�����[<N����N9e�5UVV69��
�:7�V�ˈ����,&&�2Gc�Μꏣ�=;�A% �4]��f)f�Z�O0��YN2	XkFFU?X���������7x)&���i��2&s�����G�)���Ѹ�S�[�����4��,��o=�n�6��v��à��028ص3�}�}&�A��EP�9�ab� �S��9v �Y�F#��z~������#�i�?B�c�pq�(�I!�=V���}�_n":��W���������,�,!H���κ����Q�8���"i�Ș����.�3ܒaCJE!�M���Ͻ"t���|+��KϐA# ��-@� Nޠ���o/�٭�+?������[�o	�� ������h��@����𢊂�������O���n�q���0"����>����pg"�tP�  ��s��x�����愢n66>�����_4�@�#�j`�D�Eq
��A��<���0���bq�c��nbb�p0�vv0>���,d�`��u��^�`P��.exm0/5|B�w~D �R��
���eTh��Q<f�O%%��_�E@+���p�8)��L���2˯��'�]ٖi7��������� ɒ��Ly��tQiQ{{V����111��P���6�	��[\R"
B������+4++KD��&�Kl]m��~�K��g�_N�������s8K� ���@�P��{����x����e�ץ�B�Ԛ����oב�ہF�ý�Ǐ��9=}8�<`vl�z1FH@�����(�j`M�W��DJNn�򿚐�����@!������`Z�Lv��sb�]g���\RJ
axd��lS���&����7q�/z*.�7�RRR+?�Q���,deeur��o����?�xeFEQ2V� 7'�����}�'�2�1ϴ���������g,�ss��q_�*�Nh�:a~�a��>G�Z�')������~I Lxș�(������!Q�< ".���tw����;X`E?�a�Jb�װ��y�2:1@6�r��qD��|vrq� &T��pA��9e����Zr}�����X��0�H���tbM;?��T�*E�ᔷ������*JJ�D���޿�`|�ԷS1==�P4���fٹ�����H$��y�dт���y�c-EljL�a���y�RR"YB�'+����� ��o@��<A�A,��1�M��
�1���]��L�*�j�PM��F�]�������H��X��FLث-'hP9>���F�	E�β�>����! N��fG:��f��7W��������B��)p��\���.�����A�&||�Fh((�����u8���z�6��s�����ŝ9�at��1hdBU���D/UU�0PQ���k��NNMU��}~�j�����^�q�?C�z����贉����/��D���]��&�6��n�B��rx��U��W����X��H$a���BB
�u��u�+���;��p���`���^��dd����6���VLF	�~��7W�
��0~�+&���&�ۄ���&=���;-L��j�D<�2:��&���A�K4ғ6���G �ʨ2䓐��s�wuH�9���`.�y�w��!Ej���P�>W�@)�G��'C��r@���5�l���sb���VITg������"�"�;���3:ckkkz"B0J'''+B�9���h�f*�}�x���������D��R[��e��� #U011!���.�5++��w�|*��P���Fj7��趸���m�'n%hr�c���B�->�dW��]*SZ+:C�O�m�z|�lf*t�����̎��J��k�uq�T,|x�7a����}{{{;{z��ß��z.g(��ME��S)k���ʤYA�#Xv&3�>�|0�/
>+�������	������'&�{����Qh4��T�o�c��]��i�\d6̭��F@;���##}��XW���� m���'�EDFB[O:�>��E��(iI�Rcc1��| ,���u�տ<9ɦbٳj�ʨך\�;��@J����!B�4 �B��@`�����y��+���|��0���U
?�}��������������5I�6/���bjj���3a�~��/͍�Y��� ִ��^t565�i�gk˴�;#����{X�Wc��UX�d � �D�T=�Dm����l��MIK[�؝�Yj�׷~��ENcc��0�Tw�p��}�4�����]k6���EET�>ϙ6�Â�������Z�ϋ�s�/��?�����: ಝ�������߽��I+��S�WV�bj�V��T�K"L�p*'2 b�j�L�������x���֖���Tp�O�p_]]��K�ݫoll�ZMg�R�?ʹ����;@��!��@1�[q���2�Y����L������B����Т�\81�t!_Bh������_�~�0rd\XN��}||��� &����G`�WA�>��v�����ι�D���G%"7�c5े�4���w^�����i׻���j5'Y|�h�����4�o�fZZ����:�X�nv�����v;�j��"Ds�����m����B6:s��JxswgL��BK
��m7"�ܒ���pj���k>g�z�n,��W�U�5���	B0Y�,���C)fw���H������t��4�R��:/�Q�Bnw2�X��{��w�>/�mh�X�o������W�C(|��@�������'���aX}�ܑeLy��M��@���pJP~>U}�N#�h� ּV]]�w!�w�s���B_���%`�zKT�X��=�2�-�޼Y��#�Ls��|�	�� ��Q2�1�t=���5G?�yy�S7 =�H	}*��F��:���z�����/�\_Be5�Ro����;�>w͍c&�����G'���k������a�?�����D���>���||�7���J�buBb���/pe�s�����VDG�i��Gǿy��O���yt� r���@E�`��ҸP��5�&+EVQQINM5��.�7Nh�044D�eW��v� d��x��9(=}Q1-#�����m�4�^^n.�~��$�$�����4n{ܻTZ���&�핕�O ����"��*@�V�1�f�M��Lt��~�%�6C��O�F�P��P���i�r'e^-Ņue3Yj-.�O~�̮��pGS���i/,���9��P#������^AK�����T���`b�����0��u~Ơt�>ҭ�g���qQ�6�N�HE9v'j���MU	��c���3[4�����ҳ�L���**�o�`�,l|�Z�$� ���m�&�1�Fsw�#�hhh��nQE{ZJ�tM;�(��O���e	������}E�Z<����J�\@[� PL��f3����3~0 D��(��Y_�z]ɘw�W c"�z�œ%�һ�	M|}V4	?.x-Q������b �FFFc��ڳ��F��9,�gF>�� %}enn���x�&���84$Ӿ�l��>��1 �D���@�WV�,+/?�=7��o �Dړ�-�����w��Y���w���3��88}�Z0 m����[��җ�Fti���i���U�� �` �.%�M��%�ӥj�Br'�^ q�K�w't�2���z�3��3I�B�jB�����r�-�/�0����j������������C����:����p���
"b��KWY7���5d_dt��Y�u���d���5�KlPQ��M)��[bb��B�1�2��U%��ǀXw����`��9�q�6�|�E�ut�0�!�>��Z�Z3T]���_��jB��S��͘�ǄzD�}}�����������SL|<6�MS+�p���� �x�6��NA��u<?=Y��G#��7���x��&(��2�pzQZ�E�A)y�MO&P�~�����8�F��b݇X�aaa#-YY�4.[���7A>�-ܰ9�_ccI��:��^������A�����:۲���<О!��w1��w��#�̴�m����vT��@7*1??/L4��p�]X���+�c���_h[Y���"�����L�`�����p	��� X�T�74AMDk����ᄭ2�'��H[�Y�3�_Ƞ�Q^^^��MкQ#���\T��;�bVkb>�}'�Ǔ����E��~g	����fnc�:%D�kii�8o�D*P5����e�B��.|��1�k�d.|�gOX�� ��^�x�0����,��]����ND��'z!8���6,+(��{��577^II��C��:!�Ǩ����X�
��A�,���曛�y����M1��m�E	��eы�j���0nϚ�
E��	ݻ����D���6@�=N)��כ�<�o����v�p����[�m�df~egg*�u�	|:!� �Я_�w��U0`��SR���V�f>�9R����Kd���f�+�=��`�:����xy ��F/���o�rYJ7��?R<�K�ʒ;4��_Oݼ5��98^)����sP���l<걥�u����`�+�		���:xbGb��N��U|�laC�T^_ow����^�����n�,��@��,�K7x��X ���[�Q{8_����z7B%�o`M��U�Q2��b>�&H�B���_��w�)O������!Ϩ�tq���ѭ�hii���v~�s�nfk�*..����M6���f���ƭ��{t<��+�~�c��H�
���PY�fk�����W.JK��^����@>�RM�nquu��W$k��+�����NT�!�Vo����Q�P�n�Ƣr&v\	�up�!bdff.����,|��X�K[���p"��U����'-��.�8��1e���d��mZ	1䜼j�-81�Lg�{P���\��U���̠D�טL�nצJ�������������p����ݬ�ǐ=����KR��C�ŋNN�A/��x���D%�F��$!��|���RQ�K�ֶ6�a��?E�de:M�FY������ ���c���H�/.)Y����������b�4�0EX�}d�����ⴋ���*d-���#p)�%%�����t�5�+�f;�m(�����P�y�\��J���g��do��O0�4���! �������N*[[�)���f���$$%�����C� 36�ַ(�n�Q�b�Z� J�r��(@�)E����q�Q/B�����$h��hk��l�?11[����XB@l�0�CBV�5z�����U|"v�ڠ6�#��Q��9���^��_��v|�yf���@��'>>�ag��P��D�b-v	0'��?*�������C[&4�
�pP�{��VA�����5-7/����]�D��O���<;���)"""��͍�vp=| w��B������l߷�m���76��Î����#xt����z��}z�ޖ�ٍ�
7F�1F�٥�B��#s��} ����l�Ǽ�<�����M��KQl��^�g���u���T����Ͳ�9`�"��q�[�������X�W�p�Q�ץ���������/���]�`�Y|<l�������Ֆ�]�?~pӹ)�0���т8#�y�؛B���e|�������,��%���#"r/x��o�

�^"�1C�y�����O��4iՖ�"�o�������C}�O���=[���������Ys����#���ʯ����ȥ��l{�?�lFp�>�ݎ6���16�a4	j^���C_�X��M�����̙���N��2_s0�F�bG T�:^UWIΉ��uSj��W���8��")��8��ccc�D���E���rZ��+f����	˰�"a������%ѽ��...K�,-����Yj�xYy~|pLzT��w5v���5��ڲ��k2��~
���j�����,��lའ����-&���瘘Ь,�H��X�ϑ��l	� ��w�=h` � �n�vbe���	��D<,�?�� �	A��7j�b��>ݣ���׸�綇O3i���U��a�֎"ZZ�vK���Ă��(��}���1;;~I L����GꇒDn@)�W��e���N\���ך�R��xj���႔�B����������B���[V�O��|5557�$��t+�
[�O~�$����!��WTV���Cl� 3߮�	-T,6:z<�qTӐ�w�D��[9���VU���/�h��}��\�%hu���b��b��#�.g"Q�@�@ʐV���i����<��ko�+>Ju= ?-'ve�$v��r48���0��o��		��u�i�h��l�C��t[�>�l�]�B@�$� �����X��1vm�((���]11����13�1z�i��j�^�\�yl��g��)������^�e�4�O_�W-LK�bpWy����:�\�;؆7��^�2�o�5��N�9-����*�NL�����,j~�"x[r�&J���k�\�=���`D���i�Բ��hii��4��988����[j��H��w� ��K���r%#�@M�N�<?9���8���,.��������d�3y�& ��TT�F �+t���[kj����V{¾~�zc�^1��KhWL�4/�u�P���O˹��p^�f����.�{O9�aHԫ���Cg0=��������S�&A-[��VO�\���2��|�u>���"���\�ɫ�1<�=&2*���f��{�DDC=��7)SQ[Z��=1>�ۮ�y}O�����O}&�l�C�;��]�݁E��1$��]�#�9��t0-/g*��F�3pw�ș���!D��ꃺ��{i��:����X����y��X�.��M��^a9�f��&0(��&Skf�[�$aF>Zmo�YDS�D���(�R޾��L���/C*�F�N�vm$���zٟ>M���M��C�8�K��Nl)�`���x &��Ȍ��7�����;��i�䄰� ��ss)p�޾}�����z���B�［���Ј��4l�^_���u������A���"�����x	� �XaP�
�||5�����85��n��Qg���;C��|[��r{$-��ug?h}�o����r�k�Q�%&%-��}yyy`>H�W�BG��^��եC�tyɱ"lGE��Z^S�|u���ER�t[�ԍ9��%����	���g:���`���z��2�zw+J� ���18�IЮ%�X���W;��xE>��[�3R��v�Wd��x���B��~��(%��-8��e���?C���]O1?~��������m;�6M�
����꩕��L�����BT�0�vi���zN��TZ�:���6���h�p�M�9���������w�V�SZ���t?��+9յ������cĎ��"��������h�?h�
<T$�=dST���r��"�,�[AUU�"w)�8�?1d(N2����-F�[
�2��
�~������«W��_Ȅ�����[h4��k���?�-!͋�W��]�.�����F�oko��$Mdpb�{�L��ח�j;�wAuB(29���=^ލ���K_aE�91dɢW]]�0DӦR�w�n:Z"���c�V�B!af`k$�^�i�ϟ������=�U@8my.��vڔ�Yw�Se3�����_�d�c�,�L�ۜ�T?n���g��M<���:��;<�/S?����8�X��m��E���m�:,X�қ���NwW;M^Z�3��W[�xÿ��tM��:����\�����(���F�x�՝���e��ޝ�S�.�n˳?�>#�G�3�뙾���n�%�/P�2�x�d��~������2ʬ۶�YTM)f�6�:����p�>%�� V�����H 3�֠�w�rt��s3��������������jj�P�+@�����${DDD����7R�����E�=���>NO;%%����}1Q�g�O�v�%o�uTT�:;;q�o�����|��F�ux��������F�97'����"��� �T��:��/�o҅t)�+�Ov�ݵ����
������B��<��*��??��'�o
E� ���~U<����?S���s��n�	SOk���La;5�Q]����/vKG�0��z~��N���u���p��Q\O��4�d��ㆎ�C�Ɩ�x
���+.� ���K�M)���#������N��.����m�}��gԎO-�ؗ��<j���ˏ��>����~��U���z�Qlә�:�@A��>e
z;	 JZ�Ku�!��1��D���y�m 8�V�1��Q�����v�o-�0�n�Sǟz]��� ���Z�\��d#�_x�~�\�&�I[�U���~TU��N�F�9��[ݳ���^	�t�o�/�O���	1xk �9����P�33-�h A�s;�� �n8K��<�]���2�fo>�n� "Z�دWR ������&���2��[���7� .�|��e}�	h��n�1 ā�N���p��[� IH��e������)��hc�=��z�8mi��ܳss9eee
�222�ۀf	��\�,ض��րW����,Ƭ�lp�5��-'�ru0�S�.��F�\��,��1|]� ��:���f��	��ʛ��U��~|�X����_	���,J��i���6�|�.V����qV�E��JT�UP�����|$�S ����94/�T�=Z&� ��o>~š�}WԘ�z��g@�X�-��=On��0nъ�Q��g|�zRť����XB��$Dˉ?Bf��LD����*�8z_tŐ�{\u��*W,�!v�Q'$��#?�-�"%'�ϑ�5sΑ�<d`�{w�y���X� ��#d��'�c�ޯ�+O�(��\��&�9��+��T�<�n�;����t�1�۾@��YFZZ$����'�f��� ��_^�y}D�*0��UU�P����{�R���]�9%���D\6�k}�J��H��{������b˾c���ʊ���go޼�v��^�7LTњ:��"�?��:���@��3E�9-8�t5�ۗ��������}MH)+c��(.-SQ�JLL����~��g<U�zٿ��+���K%7�+eeeY-l\\��b�F�s��u_�j�.��+�:T��j"�Lh�
�X)ho#�B����������=42���a�q}�� ����w���bO���	s}����az�lbb��+����h�X��LL�An���"�?����uY�t�~0����wa��8�F{smMl�`�ٕ�1U�j����Zs�T.(:A��92")/�
=U` ���Z���߫iiE�=�!��Po�{���{u�=R�]B= Jp��{{�'B񿓋����wa��▚���g]�.X�<($W���m�ܵ�T�-��wC�ӌg�uur6��,X ���Á�e�/p��yN7��n�3�T_ɏ���u�����5���/�}h�
�+|���CSӄ:�e��$��V��Y<i�i�Y7��ͮG5��5=�;�-���"�/������|{��A ���$�4]���B����	>�����[jj��?���&'1u+�u4Sj�M-��43�C��^|������^ZZ�r|�\��ƀ=j����ۏ�":��������>�[��|y��89�1��)<<�x��G�0�~{(C;{54Z� �0��n�X�ʒ����4�A���^��z_$��P�9czNN���(��ItOv�FF�XXX��o��:A��YH{���xr}�^C��d�x��w�Cb|����ob��X{���`�~
޹v�e��LÁ/�6\�W��!�dBf�36�;w�NZ0�n^����?�@�U��弋��?��j���}�->���4oEn.,���c�'dOOϊ4|V�B�U�r���r�F��}W��BP�߽G��|�*�c7y&��<���/�o�k�ޥ�y:�D*�?-6�����LIɪLM�]_S*�рGE������lWQQA�0�g~s�/��H���0��ǜ�R�0�cu��5;h���3�z�Zσ�A��oHh��障��Z@d��S�%�>koo�V-��������k` ,�R�曹�:ku`_kg#"#�6�>jkGJ2"�K�⌤��� V_;�L`	�<��� �ZtA
m�A{���1.NN���� ��o�z�� ��-��~�q�:o��zgfV�រ���H����x<WR�����)�!���������kaaqcٞ��|�[�І�D�>!1��Z�af����W&ڻ���Ϳ���r���?�Ư~�V�A���~|�o�&�S�juI�sd$%G���l����O�q>��!J,f�_OA����(�#��=3e��׉�:���#��ލ,���sge��U������U<R.�<�iK	A,���P�Z��a���6/Nhe.)ko�J��Ѹ?*��7��Å��&������qwqh�+��h�;���j=�����φ��:hb�����r�[ƈ~�-�B�Q����	�tC���yF����]T���������jsc0;��a��(�Ѓ�8ZE����_ �J�A�9Zj�|����������O��p�fm�RxU7�w���� k���|W�\9:z�������)�8]������C]��0��b�<=.���K�dGBF�'�y�u}@	S/HEE��'��VKI5�k���yzz̴C��܏C������v��$�oG8����D1M=�?#dr+j�Y��Y� a���h%M����deE�(Y��qg5���E�A�ڮ�3^W۞��IfHe���8�}��"+|y��o����3vyY]�6��D���ro�O��V�oϡM�v<f��W"7q��;�y/�E�?��r�Z�7��z�3���C*�����O���.���>�	�����Ͽ{YYY�����5�N�Y���֬��֌���(��ɀ�A/�<��D������{��<<���T�+f�X�Ow�)�F#��髷?a�SS�S۞r4X@��޼ss��|����D�HLS3����@�����0KOO/�gwwW��P�B:uS?0h x�3�� ��''ݷ)@����i ��������:���A����-�[4v���}G4>l333���Y�V��T�h�FD��Ů�N�O�}֟?�jj��{�������n �@�� �/n
"]]��m G���k��2�m�ڑx,�Q���#��5��ʤ��wE�e�e���z^&�?S��X���_,X�I�J��8+qFs�2z�MT����ׯ0����)r�/�`s��KZ4�{SB��m�49'C�����=��G�������>�>1�ᘽb�;�AP���(gd��~�?d*ob���f#�÷|����ӛ><�wȧq��V�g�"##ML��d�Ɣ��e��5�~u�(r�O�	��UBρ���x#pb�m�JNK���� >!!'?����B��b���)���0��SF'I<j7�}���K�䔔����8W�G^���"��)���W�o�[������f\V
egWƻp���O���
b`�0����2���I���,����;Y��I�žT>���:�
_�@-��=�H���c�i�3��&�ϒN��W�����ۼ� ��=��p��"+K��|������	^��KQ�1ٮk��c�z�*+���PG^))MM�"��w�pb����H}}}t�	�p�����+&I+@���$���	��(�عNv�Gn@�at���ҟ�á6mE�II[[&b�SZ�<�����ꁐ�|����g>�۳Bϓ���օkL�:�K�D�q�R���q�k2���#�N�!��{����o3�R�w��d�>Y*�(F��-rOo/�D����o��i�V���-6l�НÔ�B�����������=13?��x�,Ɋ��lw")i�I~fFƨmJ�8y�/��p�_��g�@_�� IHQ;ĐZ[�1.k!��D�䬓�����<!�`t,����ۃ�k�[�~��_�=��%	�4<��K�+��k������-����l��>����s/JWE幷��[�窅����*��!�Qp�d� ���T�H�<!o�?��� Pf��������~hHJTI~T���%n� ����6�#����C-ԏ&Y����[�) pED/���R1K�k|�zIE�B2�/v��#K�<>6N�j��������
��WJ\X���äq���E����eT˅%�8�L8�k���m�����
R��Z���
- �qqb<~l�ڃ��;88�XBGH�+�)f?=��Aő���Q���4U�cCsi�������<���E5�/���|�c޷g� �=��M~�gn&!�߃�N��������2��Ӹ���8�����ဗ?�����2yӒ�g��W�fS�i�e�����e��!���?���'���N��)�_�x!*F9��T� ���,�7k3����h`\J_H���v��^j�(m��=��ȴI�<e~���'t��h˜�Ŗ2���"���)��H�]���y�a޻�=^/:^��ڰ��C�2��F�wݲ��6�����܅\�swg���T}��ů�%y+�k�W�%�v���3V)1�fG�)��u�d�'/w\ڰ�����vK���È��uYW�mMe�33��Z��F+���|�/�<fQTXQ��{w�EhY�υ��gX���e�lݯ�wq�(�_e$����y������T�V���̪V1tD��%L��{Z=�[���߯����M
FnG�!ȟ��%��޲��:���3����Z�r=�_���l}X�р��!���*��ñ�q���8Zh�
�0���6)���c��<='b�)��s�",gW�_���o�X��,W#�*v�z[��4V0�
OT/�4�OHظ����m�mQw���5E@D$����C�"���j-��,-D��<d�a������H��)A�D�4�iq]����}�%� ��L]�!_"�pr���#��J�\f�+;��%B9���Xl��gCz)��3=�B���9H)�UH��IW����7�p��p���/gVE�_Ϸ���I��
����6'D(�MW���_�J�*����8V�`�=�XĀ�y��i���ͽ��_��ದ�s��_�j��MUk�O���q�N������@B"7�9����m�%��9��}��y��!��{�]���/����NȮK�fLػ��[W�2ɛ�pG��S��^�a1�U���.�va�_~�mi*o����vǛ���)�g�`�_88|�F�ezݴ�yn5�@(4��3�
s�N��Jdp�7�᲋E̋I�j�(��=u�He����_��㧥o#��Qc8���v��[d}(�w�����������E#�m�|}���d0L*>�3���g� |
�7*���߾�Q����N��e�.3���Y6	hz��r%���5�]�����ρ��j��̹$)
���h�U^|��C��$B��A���kT�3���cy�XOja?#��%s#��g��\y0���$VE`��ϒ�I�F\�]&���-cH~�_�Xk��p����}�Z)۲r�NX��~�dj��-&����kO*L���e��Î[#���Z<���:]d�C���׷k�'��*b�4��=��E=�1���6"�`������$�O�u�f��[˶����m O�3����!���a9fɱz�Y����㦧K��������˂�u�i<X?8�gUUEut�7�Ϗ����<V_4\/�����x��t�D��\��/��Ȓ�w#��~4�T�h�9uW�ƍ����{#�)!!�n�������%o�`��0+��(��r �&''?��gߛ'2j����K��C��,������A^�zs'<�"�����D���v�vRb>��`B>),�����͚�C���X��k�|�"��Z{z?iQH���W�~M�F������{]������������v����#�>Ҋ��tR�/��R}�샭�I$ȍٸ�e�d�h%E:�F��lBR�bYa�~���Q#���ym?.�X����`��}a�?/�~�ذ�k�ҏ�-.|�*3H��#T��N�m���~�����~R

�[[fI�����z�}�ϊ�V�6��4\�{��K�)U��%G�(0M�B�6�ޏgIS����qq]f��\|�-_V��A'�=v����������?�F.�Ӏu��K[N
�wVzz�����0�?/�gF&����I�1}ʩ�Z�g�pM�����L�����$p���ߨ�l���}S]�5��w�=D�,Df�����_9e��>3~X{�E,�S!h�Б�p/�Y�"dmb�Ҕ�Y��?�������P���j\��t*E)�J��QlbJ�|�QJ1��7t���_�G#�t�WSuLT��D:�ʢ$��f �([���L}eT������.�%Hp����5�;'@p���{p��aqxg���~c���ꪺ����\�*/ �i���X�g7�D���vg�Hby����P�)Ooʜӕ+Ѭ���?�)~0K�p��K����VÂ�W�I��u$�w�!h�Sz��O��g~����o}*�1qh�@=��8x�.۶i�2z̔�lck+^�����}ky��O�1(g�+�����n?����ww�=����H����FVq��>���5|L�z04�KUO�r[�i��8`ܰ���	e_5�'0oȓ�Fx��q�J�z�F�1��ƨD8h��<�@�X�9���$K(�b�la:P�ѣ��)� =(�z]���
"�,G�vK]���m��IN4�"φvIO;t�+�E`PI��,�:�I��j(� 6��J((@d����_�9-9����nr�Q��v�B (��0���o�P��}Pɰ�>tUjc��^ȕ-͓�5 �2~�9��QU��0����ݽ����}^�#-�^�ZZ����,c4�m4����]A�JS���~=Hً� ;w]���g(aSk��7F44a��Z�C�����A�߄�3��%���]�:^k���0E��p����w�0��,'1b�݆����	y����������NYS�j�u�F��y;��t��/�4�ABB�ձf��W��U��� �+:f��CU��$�C�a'b��4t���_��²���U�ߨD�a�O���̅4��t���^ �t�T����:t���@�ә�.��@�E����b��mfk�m�x�So��e^��h��U��d�ȿ��g�8�?�F�:�ɘ	~�'1��K|�`%��.Ve4�},p��z.��� )!���`K�4̸B*�/�%��	@g�P���A�|x� �F�|}�M]	�������}����^-\>4�uM��DL�<�Y2��Q����שp�?]9^�r(׮�n�[�X�PRB�e`H�ņ1��Bʒ&����D wD��1�AYҼ�x=
�=*>ƵEl�E��c{�3ϧ�J~[$�A�ȅ>��حF޿��z"�n7kq�!���(�5[��H ���O�>�ת��G��ʠ=�H(�2�l�n�_t�mYٹ�+�Q c*��U7 �J�s��nˉkl2��mJ����D�T��U^~~�ՉP�zii�����UNy��ٷ0�0~����e|��zYK�,򬗁4�w��:c�p�����w/��}�n�nA�Hpq�F����*�MO�$�RNw��x���$ttt��ဎ����H�sާM���� ��������n�8�(Y���Ճ�;~��GY���+=��KOUt�m�v_b� ��?QH{g��|��O�2���NXl�etuK�S��`2���NH$�����d���@z=��T����.#P�7�&�F~S�fv�iH��VfNw�p��y�/��1)��ZOi�������ot'�/�W\IO�`'�<$]Mۮ���pv�Τ1283[�Q�keS�.{S>����l�� :���f��*V<=n�Sz�g㿤%��&��\!��t�����E[RR"�_FE	�����-p?*�v�R��@_�]rRS��� ��t�)9�霮�/�Ar�����e��H
SP�³o~-��N�Gs�p�D��z�Y�W	f+;	ds8����AC�mtfWb��ǣ|��f��AH��Q��f|�Ŕ���$$B`s��g����@`M�L�.��B�_��` Ȝ�mɊ�'�O����$OC�p:�I��RjF�W!��*C;"Y�V���N�arycA����k����*sx�
���	r�վ��B������d��&uI���i猾�e
;��n��ğexeNxs�)O���Oz��.VQ��s�f�<d`@&u�;���H_P`�w/��S�9	��W�4�e���	���ֽ���/jG����9\v��TT��Tq%��x���'�������ɃQ�R�qi!��̤b�\�6�<������k2��R�٫g��M�|#y����訇~�ʅ���U������"��e�� �`���U�[DQ�L8X���L���0�W(���&�o3�ek����
j
��\�r�B��d���zӳ�p���E�S�_>�
���a�4��ފ������9�\|��Iؔ�ޓ�����U���d_�$/Ij�p��ڊ��px��V�A.�imvI�t>����[t,ہ�w�f�c m���i��F�r���YCJjNG�����(�/��\�)aB�œ?��5).�56Kw"�p�GI�ry�qqqU?��oϭ
�& {P�� �����^��]j����[�`��~�<	ҡ���V[3i`�ɰx=�v��#ą����͟~
�tU-B�i3�h�ﲍ�x�bФ�9�6�+4��ܗ����˘�x�GG0�W�u�R�r���cʺ<4�ҕ?�w�1$��27)���CN���N��s1�Zu���MD������1�𒢳|	J=�{.�[�v�og��X����F)�.�⟛rn�i���:SZ(�3�HH���;3�u
����9[�^�W����1��������MX��{{�P�����]��n	Nax�
tQkmc���+,��ɕ�o���e�2�a�4���)����4ήl�S�*a�_��`�ͫK�I�5��l��Ɇ�pz1��' R�J�<�q�f�����F(*^���c����iz����*���H�`Ǽ/>�`vm���䉡adD�����5�.��Ô^�=�SK��h?D���xFF���-t[�q�a#"g<��I=V�X}eZ���-۴сY<�5l�.L��g�r>�޵�$���Q�u��L��׺�A�L/E������Y�(G1䜰�������_���R!k_�R���P^�C(�h��ִܗ]��U�r/oΘ��&���abN�&Tɟy[��	##����g)�zo�A��(K�,(����D�#j�7��R����ݱ}e��oN.�<n1�,+�'fB"m�"�އ蹼�ܶ2ԉ��:u�+'N+�$����^+&�(��	-���^������^�#�[f=l��K�N�&��L�0�v�0^��y��0����X!خ����#����$#S�4{���������UsY�q�_^}D���bd��ޗYUir�7�᠈��o��i֙��b��y��n����}U�zg����	��6:�B�Ff�P=_����� c� ��3��laC�y�s1R�����K�W��1l>R���C��B�s��YQ�T�䖯����~�<6����ԩBN�$�ŀ�:{�΄�%D	#�k�l��)�u�2rL5�G��K��T���[�xb�TkN��.
��d�۲V��120��O���M���T'~�����Ƴ�zn��\���rdG��nǌ+;.-վW=�{|����'7�M<Ӑ����|��F�~��7����"3�7�ל�tx�R��HB���Cmt��rژ��dB��%:(f������[��5@��e:���N������SfSib��	�����d�Tϱ��j�	"���+��ʮfӿ����i��˂ޱGr5T��W�+��O���q�G�º��� �N>-,,���;Dd5�
~������'��m��N1�߮�
-���V�K/�:��X��Q��"�P��a'��p4�����&v�׏ ��߬f��Te3!����V�-�@���RH���y�A��9}��AǬ4��*���M�؞cv� � �����Qa��;K����8�:��"�UD(�>����O��Q���0�$_��\�Q^�5��aAWU���A���������0�҂���q������!(��km|�no�=����/s�xi(�<%�锖���H��Tu�.3gJ�J9Q��4���=�_�L���\�jӆ֠�Y��𲽉�d�$lo���/������;HWh�D����s����o���p����q�?�$R
�|����Q��E��1�kqFT;�x�RDO�o�3|A#�'��G�P��b�x}ѓ,T���҄�	���X�`�Фp����������\+M��\�ް2���Q���~���4K%~q��F�Dz�Jh~�ڒ������z��iaFÄ�VMGgF��q>����J�ٞ�8q�1��fOHޜͻ��~#Id�!;̱tn�{�#��g3Φ���+W��B,s$+�6�����{!r�!wQ�����Sg~�4>�u�>�w@�܇|��1YG��|�~�M�4�K�����[��:aI��¤�h�)�˾��Rp��(�dH�TGV�7���.
�CV�o�9.XRVrtG�f���e?�n��Sש����,�g�Ӵ�#�j?|�W���
;Lw�˭ F��|�Ϣ�9����͠�@L��_6�4WHӡ��<�)��Z^��h] h3�.�1���ڎ�YM9e�"���P�0h�PQ@Z�49z�L6O�i6��zܖ��n�����0:}*j
b�6vd�D���+s�+&��gzTS�|?`��f,rV�OnJ���<��<t�'����$bBN "I��"�@�!�k��$)�)"A|���,z9����-a�27�R��
�P���,g�=�I�Dܨ�tgf"�����1(����ǰ�����Q�{�M�__?������*r�gd�#�am�����yî���s;�֟���H�/a�C�W�-��{��M���r��d���+-ke��1u	O��mme�>�n`9��,9���FG'�[Z'�X����fO�֬$�E_�2�L�s���q���W���C8ox�]�����0׈�E-w���R�e��=)�fIa(� �Y���*GQ]�H�	g����e�_B�D�nhX>�b�ό{g˘���2j����g{��)alr���Oʂ��V�>�n����Zk�BpUKm�>ic�T}�����N��ښ�9�*�WZ�逘�'�ޓ���)�������G�x
S���x�R[+a)��L�h���37r���<	��������HCr��Q�\�;��"��ƭ�w� EN���5���Pm�l"����Fy`�l�G����k�<�O?i�.�^��?3���`����ӯDF#� hM	�@xW�$�}P��|�B���L:����ݑ��=wZF�g����hvt�+%������i���1a�l��GL]��b~��� �:�����&�Fb����|����8v#mcu䙄5+c�p��ԕc`>]APf9��Nu��;�k�>����;��!Xg:"�7�ﳻV�����A�d��[������\���* ��1�4���!y��5�Q��� ODz�_��-���'�u�E�s R���b9����MMi�:}���j���g��{��}P�dk�9zI����|���5���X�t�H��\��Tp� �Pr[�V��TV��� ����kLX�<��/u��Xl�8V�����甏W`�T�[AE���[mG:��_��� I�U&�p%,7����Nf�]؆Q1cӟKx̒��֧n�l��Ewh�Y���lz1u#4�N�x�^���%$�	��[L��D �s���u��t�}�����qu����$��aE�d;�8m��Tn�mY�j���;�������c�(jߨ]�&�|M��н��n�N�t!���#F����øq^�*L���3춰,���ͯ4Nv> �մs�����V؃!����I��%�A�u�@�
��{���L^Շ�/q��3���u��-�@��蟇v�ͩ�YSz%5��]Z�.���6{|,z)֗;hf�(�45d��EdU�,��tXsH�I+#'w>JK�[%��ccӦ�K�$��z�v�$�M�s�b8[0'bQUۤ�k�>�����LX�o�)��X���ފ��Td�����7�#�R�9��Ζ�/̏�z?!sp��M��bR �?��4�v��/�&|Z)�z
��ۋ|����0���H0J�c21�bz��<���6k� l`��8�#)F@�@�bUF6���s6u�v���R6ٱ�+3�D���Ј�]�oR<;!H{ҳt���71 ݥe����2�U���
m��[11eˑ�l��6a�p�¯��ڗ��W�͂��]�o�ʥTj̷32�s;��*�g�.�L_������}�������]���/3_�p�O�����z�W{��dj+��ʾͯ���G0K�} �Lax��|�5�}�H&�I�ݭ�HN��Yю�Z��b?C�:LB����^)���Pn����΀7�ӆƥ�뇄�l4�8�|f�\ӹ�R�D�������
۲�i��CE[�3f��I�tQ�vu*?M��i�9��(D�����'��H�$��F���8�-]��>��ފ�	cr��^JQ4�N��������[���lKKX\I�'������Ms�G���1�aBŸ��ƫ�>*�.����*՗:��"��"���3r��� ���*D~DW�W�Ս��"'!EG8k�(�d�}��՗��Q��
�^|[��`P(}]*�v�`���-\��/���ǌC�"P���*����չg�`��~�ʭ����;��k�~�L%����#���f�P�T�H������^l�����q�zm+���.�^>�r�;<�<9?�\k�sE�m���� �t���U��KM-).N�/+���<h&�~0�o�7�B��J &�>��Զ��b&^ E��u�5eܭʚq�x�w�0z�%�g|�co���q��1��4:����0��|�!�/+��̝'*�����{M{����+��Z���޿��2�% 6���V�[ҳ��䈢Y9�G%}�Ϧ_�[;���٧��T�1(��`AFYߨ����^.���*zԍV�p�|�F�I����9b�0 �QT�PP�b�]�}��E�a��Ɍ
�b����vѳ���b�s��b��~<��	7{���4^�p�o�g��%����v�_����'s��`j�LU.�@�ȠjWw�f!�-�?Gi�<`��zs	5�w�|�;�p"�M����g�>�+�g��Č��l��y̓�D�C�@g�t\r��̜�uLL\�>u�32bj�D�\� C��t0G�I�"��R��є*�r?d�Mvq��
��CJ�@
?�����e�#gaMs�D}��ZI���x� k�!���v��������ḯ�m���0�O�z�@��͉lM�ڦ$l�T�в����gӼ]���hsk��2��~܀����8�Q�'��V�~m�*J������͋�Cc7��5�n�z��P���q&5�1D0��Үa��=~ Ϻ>�ÿtM(�Y�f\�f�8b�ohZŰ��Vk[Nc�.��(��BC�R��ZAɵ�#���}�۫� �jy+J@Y��?���9�*�k0QmP�^ �׳�"�t�*/�w�!��;9x3�]Йkoq�QR��-ɏ��d�� �OJJ�ˆ��ӕW|�Y�������O�E"��U���+�0N�Q�`�FϹ�V9:j���GAT���O����Cn&ٍ�,6�P�À�~Z���E';=6�3N�u/���!]K�z��(&�����5�[_��u�pg�잂vXA� !�ɫ�*��ǀ��E^p��j�	��N��f�!4r>���-'	kiIsӯ�U��L"bŧ�m�|�nI O��;ҳ�(j�d)S�4���A��@�Yτ �a_/�Y<�I����kZ��O�P�+����@���䌌c/�6�щ�|`�������H|���r��0����v��ͩ��^����Q���'��e�p����{�)K$�|~�y����<Ң��u�po�up[*�:_J�b���NAs���m���'4�S�;��`�:��={����
�Ikw7���8�ff`(�k���:��'u��/������`ݥ������L
-Uχ�3r�Ɓ_�Fi�Щ��,YIh=LvoS�Ӷ".7�
oϓq���?]�x����=��e냶�`�S��Å��C[G(@h�w�{�a��~��B���k��H����ˌh#l.c�cv'�n'퀭��PW���Z�i�ri*֊�Q����5�iȨ���ב${d5�[ӎN����)*5�� tf�NO�y-��q��>Yv���x�����nl�}��(����0�@���:3��e��Rɀ�����73�5���ݽ Ӿ�|�YvZx�L/�U��>��4P��T���%#$�	o�{;K�f�ȆGG��>�C���Q<>�j��J�q��L�Dn�*�|Y�i�[�����1&٩��v"�S3�{��=k��O� �=iٲ}��|���I�~����π͏���0I'��z�z>���W�J��/x�3��Յ��u�4��[W,�Ya"�;��Q")�J�O]9@�w��=��)	ƙ
c?������� �k(�'N��� ith�嫏�(��*�L藰=�Vsz^�q(��Q6�^Â�
/��bo�}�Ҳǭ&mpC�%p�O��m�r�3��U��l���/v�'@Te?���&��U��o�p�&9���/��='��٥���_4KP���1H���U�S�������A��c�^��l���	o�ǉ�����OYV��߁pqq;��.^d����gܶ��<��/�\��d}ܺڐ��Rw�����oN��D�ob���-���]��GK�
�I���	9{9�ւ'�@�t��d�7+�GɛI�1�M�Zv� PBZ�3�G\<</7Qf����h"�:1C2.�,Y����S2�)��`f��2�x^�`��3���)_U��,��%�==�O�*<�G�젓�[I�]�����}W�jo���6l/�2�
5z�4�Lk�?����_<1��%��m��Tax��氼�ϭb
@;CO���;qq����U��؟:��e4 �����)������T<zu�~�o�e�D(h��"ʟ�3$���2�Ma���_�jx�����;�u|}�"����N�L԰2�tTw!Iu&Xa�O�;��ϙ�
WW��G��m+����f�|vƔ=�iN�R��=C`HO���8>:�+�}�v�E|,O

�o$�x�y6��V��F��獽�a��C@��;ã��|,t�/����#��ٙCIY�W/}rT�����V>;~�os�zt�v��&,�D�%�V�����9�.󌀟���8L���;�7��u�4�?�p#�o���P���E]-1�M]�IQ�Z.����{g̙y�Q��X��[�Ŀ���r��_����A6�M�>�δ#�Ulc��2>A0:��������ל]#�d*�>�D#��/��+m>7���xuι����W�(�i���='5��ؤ�;?��ϦuU��2j�V.�����E��ŷ�Dw�EI��bC�U�~�~ #��7S<������Œ|h��Ґ"���}a�&#�v`��M���Dև��:���ߏ3��ll_l����N���_��M�$��9�v�}[���3]ĳ��x&��9��!�;r��Yu.��
�t=�&i1����[��~�����[Ro�ŀ{��
6��`�Ұ/5��G��d�����s�C~�s�4K�!�I-qT�&����"`?ڸ����b�r�3^װ��^	,;��r�i<~�W-��
��e8�g�V�gS햜O(�*E7e2��Q1��N�L�25x�dDO��.�^7�(%���]L2D)�u�CN�i�-\�
��ld���x���8�=���/p$en�:J�v�4N�b�4���0}F^_�J��F�����ݯ�v��FӪ~�[�����HX	��K1�<5��]䂟�Uq���5��x!/ro�Ւߒ��F�&G+����QT�-l����k3��`{<8�r[�i�tU��gN�ڻKN�Ǎ�Snޏ�������QH}Š��]�t��U��:k��Z|���m���d%]C��SڷEy�oϑAj9��}���v��p�����^�?Ϻs��U;pt��1�`�nI�M����:��9������ti-�j��k;4��A���������,�=!@B�[{����5ьd���b���,X�P�����8��H�q{/��(�*�&�t�+����������M_���A�|&�2;Zj�=�@VI�8u�cu�M�:gJA��Ng��P�-.!�ر�tR��)� �q[�V�<��\��g�f0���=*��G�����5��8Wv����V+�{CP� ��7����5>�!9��A������H���S'?�Ѓ9���2�����s��CU0�[���g�d�px��a�Mz�Ž?����V�3�h�U_�pD)�J�����{�>aMV���RǉAǈF�N�M���G�+�:]�1�(�g���?��U`��������B3�(��=`�ȯ��fX맲%o�le4�s�����Y_�ϙ�>��*6q�%���sx�'8�Ŗ���p��wg� ���Ʒz7yo!�a:F}J�Y�_/�2I;7-W��`��7D�44]�u�5D��������H�}zb��H�%�xO�Gf�VT�R�u3��T�ߵ�*��m��~�NDd���F��#.%+G;k�*Ԑܣ���<�1G�W�d[���Cu�I�̈́�܁ܭMf̉|tTͽ��pÉ�/e+ȼ}��E�͊���Bڙ�7zx����(ZC^����ps�ϦEPp�6N�Q�mq{h�j�v���p�Z�gn�W]�wě�=?z�>��1<�E�!]��ȼ���x���,�#.�l޴�tٿt./��l������zؐǣ,,	��]����<����:����B<���X!��+��4���=F��$���5�������8�>�:���Zr��:�'�.����|�YS���H}�Cq��$��U@�b����WB_������`�e��������>ZA��4Vs>�����jE�m#H QH��:�/��u��ƫ'"c�x���x�C^j̤����d�&���I���yߺ����bb�~}� d�h�,�kݛ�U`��Nۛ�������A���%�4)C�z��k�E��O�v~�\a����f�U�@�݁�	Vs�̧e�D�s&F%`[�Z���:���pi�l|����gA���f`�F<gZ
�6���\9qʬ��+[����1�V��a!h���1�}��֦VV���aadg�-����=k��,"X���a�Uk�L��+����ĸSH9Z+�/�xLe�gc�0�3S
��A��<�_[�(����ER��ƒ�x?x7n]�����;FF���>��I���>�2lQ�J#Ԇ�r�2ʪ&w���s"��K@�a�o�+�fEYo�&&I�^��9�F�R�A�J�	iR*A���V�&�Oǿ�x��I���\��rٝ�����Ku�v���n]2sl�"l��}��O�$�e�V��ፍV�����>����B�-3��
��a��­�XFjs���m�(�t����$2)����U`=��(��ٳ�Үs!L�zF��U6����RT�V��t�Tz@�[K�W�l�'��L�͜��~�	Mz͚m�O��&+��0�VS��?��}�I&4k�����u��_c�r9��j;�W��#q��5a���}�S�2��C׃�ߣ�]'~��N�s��R}��w���{����J�u��cvv�U� k�-c��4S��iՈo�V72:ƝN���la�	wꯁ	J+��K����}�{��G�T���`t{���f2�hs>�ܳ���N�v��1�8����{��yc�:�ߓeH��i@��m��ނh��Ѥ��~Bvu�掆3�[뿸����4��J�%i�l�d��{)�w�Jlt��t�vQ$���H�[� D�8�^����	%c�&~%;):�z�U��t)�B�r.18���w�na��(L�zl��_��*��?'J�)��(��\�HW:�����w�V��I]���g;_�5�L��G��O�i�Hk��%R�W���223߭��(fA��ĤD���x��r����'M�[;Lk�s�Ln��S|���^�:�����v� ��5����:�B��A�ŸX$�R����\����`
�۝}�Ń��9+>_�=����`�c����A�K��Te�%g�������(6�@����Tך��o}�+�H�� �F)�^����2:ڝ��nCõ��g�w���xk�<1f�T}_Y��c�}Ņ��$�H���#)����6�g39ZDX��?#?�9c��е��h�,M{�ǥd56n�=Ls������ʠ5>�vR��zD��x��6dx�����M�%�!��y�R|����|o��p2���������G�6�U��������x�5WL��О�9b�od�O�n3�&���4 o~zJ擥.��q�Y$��ICQ��J
��ñ7���C~@O�W��~3�%Ŀb����S_(��F����D��m!��m�"6��K/*�XP[L�C���@\��JP���]r­ؠ������w�Xq�dCf\	r���w/�����JX��c
PZ�Z��<��7��}�ToV!���[҅�����A��m�Nr�,��_QE�GX��OG]�7����TOx�KbZw[����-��'5���/1��tyw���?=�luG�������*=�@��'تj{
J��ҍ���=�5�*�z��p?Y��}�c����2�$��S��Z��)���P��H�R|���1�@�#o�
l����EsT�]Z_�7δ�, �|��WP{g6n>O�ݺ�3���<:.ƣi�{3Up�g]��;�=������uK�G	�L���޻JLXP�Ǐ�eeѵ		��d���R�����gr��R_&�q�yX���?�ϮO?QІ��i����F,��Y3o$��r=��s3v\_PuQ��� �S���ᆸIU%����q��C0����.Ĩ�� ���������!��/u)�e�RY��9�ņ����/�.n?z	p��Ɏ=H�������my�r����=��5
M@Ab q�ٕ�f�@j��Ɯ��T?�*��'E���|����ٹ+�����z�ؤmgt��/�f���fR����x]�a�ܢ�;�&���S{Ru\W,�>����P1.�g���s�o��K/ӷ%��;&��u'ߐ�X�w���e~����+h�f��bQ�����Em�RP�̇�Kk��˝����D�>�>����V���(�UT!�-�\	�&���:��~����d�:������\�x��V6g�V�Z�B�N�=w��|�DA�˹�p���Hǉ�)��,���Us<�{�/
<��n�
m$'�ڳ�+�W����ʣJPcI�b�L��5>?3��qp�����<4�!}6�RMF&����xogwhw���ķ�"9�?1a�`x��@=K%.O���:7�l�~��vt4=�~E�%����[̥��AIW�M-|���)WyC֧�9O�991^W����v*��T|���(E�f6I�N '8��́��=�8FZ ΃׆]Q�#�Sc453�sE|F6�)��R��U�a���ڢ{���ݝ)��^z횇����M6���n9�����캲{�I�p��\�;ɻ޻�����z>s�J�#�����*��`���w��=ٗ��[�a:ʤm�ƒ?��ڑ8�����ʓwD_�T+�;:dhOߧ�4�}s�̷���q���{�9C�|�$�/����͊�;
���?�X=��Ҷ�F����~�`�Vt����T�U�G����e+JI`�R�+��q��ő���g���#��oƼ:��<8-d����_*���n>���)��Y��͜Ҙ�O�}�_
�;����������xa��]��jT�����Ib���@�u���I��p��pk�HAp
WpsV\:q4�=��o�ja�{&����{�Kf��LҌo����n`���
׭�:��׬����y�n�c�I����>@�IC��$�N/�fO6�:��r�L����N�Gf���������=d�]0~�a�ѝڡIݳ�`��>3^��?&�v�y��:'�	��IK���[�xC�c�cq��#o.P�X��ղ��N��Pg��4>�

6!s�*'�����I�C�_����p�'5��3�캹�e+��q��y)P��_�$�o3c�&gD����_����Q%	�6T��"�`A�v�����n��R�e%�g�U�m���6��X���d�	k��m8HSG�k_AI�[|��*J/�0{"
�G��\D-������-6p_5hʶ�Kv�������S�2(���~?�L���5fA�������4Ӱ��%�s���duh�H�]�1|9��B�}g�]����xz��ϻ3Md�����[�R�e{_�O���I�Ĕxg7]�� ��nvQm/zf�6���y%�@y�~��9���D����2�Qݍ^2q{\�%Y�4[Cݍ2����f@�$Sꬖ��*^2����P>3�׷�1��\:�z0�X.Ua��n,g�,{n��
D<��\$u�-u���2*~텕r*F̖�p:�_ʆ�р��ުp��}�f�f��M� 
2��՝uq�LP"e�1�Lèb��@�B�#i��ǯ���q���u�y%Nw�Ps�[�K �ߚ�=@R&���B�=�4,���m����ބ��#��~\�2%��[ȤI��S��ٓ6X��Y��n��
��ޞ��^b�spR�+*,��%��B.��/�5WpR��%�����
��\U�Y�;@X?��n�9FIS�]��Qvp�4|]g��ui��j���-I��(��>�v�����������NJߍ���%w�s�싅翲���*�WM���{=�A �%��%\��� w�t���xR���gQ�uԲ#Pc�`�"�.֍�;���`�V��['`������p�0 �iϫgЇ)s�=zlǣe���>0y�ډ�%�q	�R���T�и�"Z��F��N`"|i�	��H��	U��G����z��&"���1���E�^Oc�+/0��A�9_�5\�S��n�C�΅�ڢ�������.Oƛ�d�7+����;��H���y����+�*�}ro�N�Nzo�N���lX�H9[.<�<�B$�OO]b��<��e '���m���֡��^����a���=���%$�.��h�5�2��{�v"�:,"`"��A&v��T������ �"�**����3*�c�o�'[A\!�l\���a �\P�$_0N�M6f�*(�1α�G���/�m�ap�!�/z����g��ˈ?i���ʙDb �=l|d�/@������������)�ꎝh%��V��Gъ�+ ��4XH��,�:)�󰐥g u�T�=q�~#"����G�^=�+��`��h�w�bcxcyk��xѵ��� \H	�����R�Ɓ���c��>3."�Q9:R��z�u�j�g'�k��Yt����-���lPX�0��y�I�)ło��������)D^�t藸n@�ݦ�D�i����;Ƽ�>�|3e������M3��S򶭐���V��qx��R���~�?�M�h!��S~M���N���[]I��?��W��eI5)E�A���#�WA}�O\��岆^����������@ �1�0�N�2I�c��Xy����q����ͳC>W�(�%��U� ���׈W����eslUD1��	f�T��$/"�X�,�����*[k4oMY_7����+�Ο��|�;d��J�"�E�q�"���|޽���\܄���r�4�X�L�:������Oի�pwN���xo��9�5�����5e����"�$����&��1/�F�����+��#�R���*�m���� ��._�>�%R��=;�OQC�AU�o��)����v+H$��<��^�����oh���x�m�d���{4}�`�9��
ĸ[�����l1���0ᓾ���_Wf}}�4A�2�V����oqȟ�tG��h~R�ֿe/��l"�t��z?�Q�����c�z>�Mz��S��hm� ���٭U���M������|��QK��/�O������3ra�
��S�0�)���`#�@�	�����>ӌ���D�/�	��O��=Q�Pp�՗|.�J��Ȳ�,�JǺ!}^����_��������6M��2GN藋P��B�	�����!h�'��}��G+���:ZU�.���ZedOf^e߸���*;��0��9q�$���O��m�K�̼
Z�l���& ?t�\�	�6ܾ<�k�����l~�@���	�6k \�� =�f�8�KK�Ϟ�L=�f��tM�6�2�w_@���{�c) L�2����*A�^;s`Ѭ�d��ƇX�{'{�+}��\׏,��<bի�]�����I�4Y8��me��a3��!iX��]�qbm������҉$6e��&rH�[M��#J��,M��=�#���`�*��Z�P��xy|HC��ay�`9�B�H�g0��ި@�G�?��2*�`K @���.�{��Cpww����������}����Ιs���[�~R]LO~�]��O�9:9��cA�bw� ���	�����;$�2-P�T��Qʕ�z�{��?GI	h~��<�A!�9)lK�ũ��L��5@`��+�����X_F�p����,�N��sq�z5�\�J��KaU���Gm.�`��In�A�8��pF��7;�g�DȊ����O-�5�ƍU�R�������_Xd&��FAHd��\����7�f �'�qTmoq���EdHr3�O���"��j���~5�W���W[b�uA�o����X<V�ΐ�;����c���ɔ]�5����9h:��%3ӑR*Dt;Zp��|�SZbfRbJ�	FMA<]Z+�������#3����=���C����X'북��Ƴ-����s��Q�:��I�����\;zA~�K�O~Ge�v%��6�+�oY�;%-uQ塃`���w7[�?K���3�F	/����9�p�?c�Y	]�|P����		�6�s�q�X`�ʥ��2�mn�vE���0r�nUJ1�j�����b�=�#����3����XEV�*�����̏�����g��J��ppQф�����w��^p�RGh�%k�q�eED8��HT�z#a^��.�+R��]�>� Is:M4\2�+��FQژ|��xnà#����E|"���i�,��{7l�	*t{�V�Hd�?P��)��7��/��\��o�hΖ] ���`����FGFF^պ8��qH�W����?h2��6�7��d�rUH�b�~ZiHK���Mv���uqQ�0�¤���º����o�k����^Ͼ��P0��Q�jo�6JL`� �I����!���_^^N-������DE�
5��dL4$PCG��Ɇ�K���9YE(K2M����KZu���;r���兖�c�����!}~] �1E�2M�
����-�?'3�>l�r~�D,��k��۩���B�OJt�
�>pV�	���6'trEƟC�����Ft@���H������|�Ԙ���kM��yNNYY�IK�׍l�A�N >a�<��[ �w�;�c�'/���:p�81�|,�?J�;<R�R0��a��C�ڟk��
��
����[bazD���1b�B1tA�k��>���B$?�/;�>O�:�K^ b��9������#�z��� �&dF	p�ρ_(d,�?;��(h�}l�\J,�\2?Wg�<�+Td�P6�l#�D�=`��<Cޘ��ůP��/��Df�pu5�m��3c12�Ŏ�4ڞ4��￵Cz��F�o���!^r�)�~�5Yocq�}=Q�3�@P��:�0��i3FǽA$|���y�#q u���ߩA��Ki#Ռ�ъ�Y�N�C�m"G%4������#V��B3��Xȫ����ݐ_m����e\�k�����.�<˩y~O:CJ���t@+ޓ��%l�m
�*S~BΏ�d�=B�/	#� |��x~�%�3D�H;�1��N\W@`�@�_M���"c$ˌ���ͥa�`q��iS�Ɨ����_�QQ�2���j�3�iQ�>�c�|q?�h�`mh^�E��GDC^B_�|ɻTK���.&�>T��D���uF.�-s��bKU�
`}e��8f���W`<���[,��'�rj4�I�iw�%w�0�lj�
�U�<)H��`�U��-�C����Td�1sC8y���\�7�\�31е��D ����Օtt�!K;���w�6��qc�V���oKAG���Tm�(�x�s�%`�Q����3:�Z�?)�*��[���]2��a"��LaB╆�E�e��s����r���c0��ܣ� ����`�@D�A1UsT��f+�c�����l��7�R0=j��Ik�:����fl�<��ǂ|�|EQR��Q����G
���%+x󱱨�+:�! �tP�$�;���t��E���B_��EƖ�*U>�5ط���o�Z�~FEE����d ?�2d(��<�2��Ř�N��Ūۅp��ћ_�Ȉ�������g���t��P�p��D�8�WX=���S�ڱ����=�bɣ\�\�<���޴����ۋ��Y��Zx9�zҤ���]����U޺:qk:��1:���3I�8�7�{�Q���ϔ7��!�O58�m,��V�N�{C�K�7��צ)#f$�Z(3Y�\�m���M���-�P�\��\QI�:l�H�mj���Dňn�����R�2=�-�Ov�,�����X�h�\����j�����PS��0ot����	7����o�f�Kk@���8���;<�<��`t{>�T[�)u�x}m'5���#����j3#v�!�y�wb���VA�s��ž*Hl�Sf[�3�����G�r�nYMbI���5tA���`��a���� �S��(ݱ��g�u�{  ֌=�ɒF1�}��hR�i��?��Je8{��r�j��?��|y�9D�Td*��a	J�Nc� hc,/����̻�zxy	x�1�+�	:���a`b �>}LS��g�g+AW/��_�_;
�k=�B�	n�m�N��L0䦏�'{b[[��������_UdU#�i��ؘB�0�ȺB��ZYM�u�uJN���L;�`(\���/T��.vM�r��:�	�I�ǆ���䜺�9���w^OܚW�w'գt�Q�w�)==5'M���e�H���vu��y����J��aJo�?(L���{`{d椢$�=��q�2�#7;�(����@�t���m�h�?��R����7�d�R��S��fs��+����a��_� ���s�6{1��A �4Ϯ�k�Fѕ�1�%!ZZ=�i��I�κ(�{tS�H�k�S�k�VDP�*��8��A�c����x%ẑ�$>C*�����N��T���7~T"Ҕ�r
N�r�@˙�Y<�1"[ \5�[,[�T�sn����`��q�6<�m�aaaQ�1*�Z����C9�
'���v��F��{�%Z�����.���V3�� ��,L�s�f����a��ꪲ!r�!g�+��
W%�E�-Ϗ�����]��mZ�`�L�A�3��3؅����zB�t����ty��^
�M�VS@��/�:~m����#���_SPG��3���R͘?�L��1[�\w}�܄����P��ӳ�����!vg�Ĝ���_0�$0�UX�W��ǐG!n��*O�匚��fv�/T�"n�[(pk�}��a�6�����i)�u����Qϛ��YA8�pW ����}�u,�(FU#���qe-=&�&����2<�y�����1'F`�����o�S���6oFo	�	de�o7�2b�N��wK(�nF��uOD>PA�% nq�{�Ay��t�H�D�X��ć�\RI1տ��'0<n�=_o�<����z!�����ܦ��1��e㜽X�=�T�(2���Tp#@����$ea��v�&����s36+�B��$�~�i�T�q��N�D���R��VVb%�K`�p=���R�W���o��Q�T#2���/��E��땐�-}�^Tl2r��~��]V"�ٿ����dr&�]Ǥ�s{���j��C�Fug./y&��q��Ym�~������X[H�PrS�KH����W�f=��E�=��H�q-		+�>)}T�����"l�%ߥ���7�5�Xʨ4��f�H���,�]@9��EM�<���NMeD�W��DΕ�66����0;P'�-+YC��b�L����a�_�J��:�D�pJH촯u�ɳ��h��N���%~����UPWVU���ｘ�wiN��A)i�`]7��:Ҧ�՗�d+��-�D�/J�]�Ƶ����/D�����Z�?^�v�/W*(��i����u�N �]Cu ��>D��j�}��@�{vRⶭ�uQ�Q�7��.r�v��wbh���^�q��@ފ���ȇ^�&:�ټ�KO5�q�~�����^��!|��kq�L��-�$f(/L�~�������p��e5�`��/dN�XA��쨐�u;� �/�dr�%\L*�c+7��ξ�a��I�,�;		�$^������Z�#�݅6�SB.�Qѿ�`�Aۺ����g�f_�E�Ǘ���]~�ҿ��G�!N��4%'T�x��w^��czfF� }����)�lRbۖc����sb����i�Z_}���u��t�fu�Sjw>��,\0L[EO�؈<�=�=�bK�ub%#�����T��>��F���;������q"<�t�c��ś*��DP�`$aa�m�8�����h�,=��u^�7��,�_i���P�$�M}}��0��'T��i��A��t�v��#/f�!�_^F�fr>J,-4Q����'�^h����h�p�H[`�m���wAA_�>/&�_�f�V:�%�f8���@Y�e�\�)�}�� �Ϟ��iK�Ѯ��t$g_˛8��bf٨��Wٕsh	�e�����ѕ7�e���0�����J�45"((�cdN"�s1�v�/�������;�R�k:bQ���sxnNqk�l����m%�|4,~4���2G�5�ߑĈ���GB��JpCCE�,
��	��!�Ϩ�ڔ2�,�χ�˛m0��l�����V={Vm��NP��Y�y{�߿2�ʂ�����Iц&f	�r�����/�`p�M�O���E4�ɶG��/�x	�����[b��l��ر�uڎ���o��د��`������ٲ�y2:��}]�\��ˍA��Q�knr1�!�	~d��������4_؀BV"�0��BB=�61����X�������cz�ls�ֶ��m͎�5���H?����q1�$:q��ۛB�si�O�>nZ�ϫ)*�u.
��&�e�qi�^��Q�s�_��َ�ڸ�2���dc"���l��t���`��8jt��P��Fb[.л�-
���E�Ш��GVe�����o���t*�����1�0׾05��r\�&Y�P13�z�at�ϕ�-��ˠ�.ovG�AQ�cc`��p+��Ɇ��˽Ű^���a��+������9�'�I� #2��;���hbQ������:C�}͸���͙t�G�tw���L���4ո)�n�I,��RY�׳��eY0��,�����lx�r�kH�g�W9��\kО��'�jK��ԈT��q�B�3�0��d�)��?���f�W9����N4w�+���Խ�fש,�}�x	�ZooT�E�$�Z�vQN�Ef��J�g��o�_}�������%9�M"�3��Kk�V;�!ﮪ*G��﹈�t��^��	t�����ü)~�|yz:7Ml}�PU�&m"��R"�������F�Шd)��y\NG8];�p�����p�Ǔ�
i7\s.M]����4߄�w�����s��'�g0Ϩ>���(��J:���iN���WWu/"�Ӓ5� �d�&w���� ���/���|����8f�cp\�"s�[�`�z"���7///����>�&tT�,��"t�/D�HL���E���y�H\�z�����$((��p0[T����R�ψ��ӑV&�Ւ��v�AK[�>Cm�8P����Q$�����6�4d�S���i��
t�<Q��!9����q�p��cýzzƵz��زTFEQ���2{��T��)����MUS��������ʟ[��������߀�N������Vn<�V.�{���9���������F-^�dV���n�Ki���{���Ae4�$�������Θ�Q���OzX�C[�v-�q�t)�����f^��V�C1���p���>2*/�6~�k ����2SkP{*��g�����1�4�&��h��"����ͮ��^�0`Y����v}�5>��y+���9A�Z��<p94�����3:X���1F1�܂66
i�����m���+�	ʳq������9qX�Y��J�'!�a�LF��J��d�S�OD	#H�G3�����W�_e�/���혲�E���J���N_T{���r&F����ϳ��lV�
�j!�`ƹ��1 P������/�;ܱm���00C��جA;�S�����#���ſ\eh���N\�k8"��6zk����*���i�����Wg��3v�%��U/����z����O\SƘ����ߏ?98�$��,;���^��mm���)�wW�iZ�=qf��Rr���QK�����!z|at=�t�	��=���<zX)�Zj
����ןH��ʴ���FM�����QK=��>qAp�+��e�u���R�|�Z��ją�\��o�X������a�X�ٰm*��z����f2��|�or�8�.��X�(�ZÑ켟5�����1�������A��7�M_�XyF`�� �vǝS儥�q���z����pI��$B�1%����gqGM�Q���c�g��3`,�����m ;c�[�����^
 Z��:��`$���DHg��P����拈��I�6s��&���d7/��3/ǝ}�;��R����ٍ��ō󵤨�,�z�[}�����J}��$/X���EW]ψutL�|tRŦ-�-&`��dvu�x2O3����#1%%'k�ϋ�/o����?��f�H�5��u�az�C�;�<�#"*��y`�pj� *�O7nx�TV[�	ϵ����v��blb�#C���9��k}ՇLZ5��.���26��>�f>nw�]���J+�cK:�9��-W��-�����wg�������`;g�P��;K��!�h�h,�E�s&I���ԠM��( c��l`da��cfCglZS���w��,O�7\L��_/4!^�r�GdD�@ %"�P����)�j�%���'�-�4�M�~#{�������
��f&:�̌�aO� }BL��$��h�q�������Q�X�
����m g0g�Ċ�����&E�v�ƀ�g�ȁf��:fll�n���fC܅n������G�E��s\L�Jy	dX�U�6����vJVbflij�� �{�ƨZ�Acۤ!��]5p������R� 1�
���L��A�"� u{�W�EA���(�h�"��_[��Z�)��آh����>:9��t��G�S��BʘX�1�S��9%�({)-���\#�hE�$���D���|^^�w�:����f-L-P����Xi/fw��l��6:�G{������3�����F������ÿ��c�\e��?��ٓ>��\>�e�cy�;��UB�G���G�zR�������f�6D,1q�E����_!�5�2S2c�.n��/͖�KK���?ð���P��	wm9ٛ^U˥���`�9��C�>��)<{��6����Y��k��۱�Z�8R`8�L��v��� ��q�&���-!�ǉ��b3쪃*,��� )�,o*T�Q ��H!Y�x�ԋbMQv5~A{D޷zX�^!�A$�dz# �>#��i�����3BMQn):t�Z���?���� ��&��n�1#P([�ɩ��VT���5���T7��TW���L�0�w���Z=�$i���)S~� �;��*=��&#��<E�O�8���E���͛"������Mx >����-=3�3�����R[5���̚%����i����v�<�r0������>J���2h�I�r�&������7�{P!���U��i����A����w5���+�}��P�Xh>�����!!"�=y&�i+��a_h�����d�����B��Svkq5:Һ�=��k�Giu��E֚o�~%�L��� M?�����F���q��X�"*��p�Qە�����y������9�8t�>h�)��ޖ�Z�T����$*"B�1����D�PǵvP�4j���>�џ0��&�y������+�&|�
efו6O<��]ʺ�՘[��H��_\�*�3�}bK�c=�
���V���;�<���+u�y�5����]��ղ��A�8��4��w�_��HkҠ����Qxg��{4Br��D�[>����z?~7�����Z���rT�m���}��>c�]�XrT�����-����-{�6���WL�E�C����! Z<4��d�_����#{�N��BHĵ���+���c��h'��Cp�,oYI�/w��ʲ� � ��� ��U]���� �=7���4���cQ]���y��S6�f��	p�/z־OZ�@*���VxxxP��;ψ���P�[�ͮ�W�:�G��A}�zy�e�Ǵ�$%�6E�9o�g��e1��G��4��u4�Ū��f��bW3�v�fm�J�e]t�H%��?Aǫ�4O�5\�QU��ۉ=Wm�����x^��e�q���><��W��.a���W3�v%TX�|Q��`D�n[��!����Wr���"�6=�I�6r� ��:P5զǒ�Y����F�ws{�Զ25��iet��g�M�P���^��������՜Y<;���O��y��K���9���^ �bu�~���*������D"��6_uE��l�4//7�}��%+�e�ǫ/j�������I��ܟ&��>]H=��C3.~n;������e��ʻ���k��q
z7�L������m��3Ac+�'���:$���"'/�J��x�V�eL�Ã�|�Hw�Gv�����ma����V䈗���t��Ǭ�4��% IR�^)��Fv��0������k���i�@�ܖ=��7A!!r�Ii���J�T��?��h�u��>��Y�/��;k�
�� �'�'(K
���!{�����L�oJ��=^0E����@
V^��ue��W>��N��+1�[�4?��O}Y���ȴ�_��%��������Lߝ���V�o8[bĒ@!-�pO=�x�)���3����8��� tP�r�i�e���� �oo�J"�&z�o眖K�L�n��U������"��s5���Z(;�W�.���=ws�`"C�$��:8-1yl�^��j��\�c<,n�K������7=bG#e�X.����|w�&��kG��*�g?������wJ��~H(IQ8��"ij�߃�#jJ}�|��Q��(m�KyT��(r櫎!��^�m�O�-��}�3�]�C=km��3K�k&h;����g���f��~;WASN=��Q`���LZ�7�ض�>��ЮTZFj���5A���g)HSF����ѝ'_2E��3))ipLq_��1��鲆�����ws3'�Q�����qqq��X����1��o�v}�?�.���m��+�_49r1�4��w���k����p)����b�:��u?w���w��/8�\>��}���r����R��L�b6_� E6D�c�R�	�R��,�?�����yl�
bu�t�����l�+�����т%O'�5�#/6���Y~9E�-ܞ���E�q����F��Z��=��?<|���c����=���j�C=c�v}�W�����o�§�q5�N��O$,"�=�̹�`�m��^J+�*��}B�mB�?%nϼ����&����q����p�Z���=Ua�)Wdx����k�|#2��=<t�΀��s�C��|%��+r��j�wa�+��6��'����e��;H��q5i!"�^Q��"��bɛ[Tf֝��ۂl�p��5;s�����/=�a�N�j� ���m��c��\'}Br��W5��
V\E���J)��M�������7�,��nr��8p;s:֤�Dp���CG�x�.�m���sCz���J������V��QWݎ��3��l���6����ӵU��<<��U��G�<|�2����'v��7j��T#ѬU��9�^��qy�LL»�)���t��Yw��]ݛ�),ebA�g�ɞ]�%>bz��-f�}�*�^s�ۡ�A��{���%�,���+�M8����]]���]����8��ֽm��[mQ*OZ���K%5�	�''�W��j ��9e�vO���gY����2�ܺ�x�8":��Ő��g�-��b���ڵI1U%ެxDV�� ���!h�Z�\Z[Z�"�J�A��u���sz���JeA��j��K�8�p��V��0�N�����0����#[<�8���)*�mjo�����t�ƚ�����͌m�H�)�n�X��x����S�0�h��
y���Bex��י5#e�|f�|�%z�[qe#l�G�*�|��q���~ 1���UE&x��[�����P��IQ��Αt�T��������� �����{�.u�Qs��8�؁�^RRҵ����~5um�卣�S�0JM< ���\%+��j�vϡ71��i?h�xqMAG��$~�rĆc�����;<9!���vƏ$��qqdw�K�_�\ ��zҷ���F�~-0*Ķz����N��5((��RK+�������i�C���瓊���҈��� ʝ���L�g�q�[�W���۬�����R?�s�$�	�Di2����_�#R�ȸ��
srP`�T��b:F`4��-�c�r�����n���|n� sn^�Z�ZZ��[�[!I�H��}��h�S�#W�|�[{yXy�ڈꔀ˼*xv��*58�4=M�_�ids6����Gӵ���\��B::�������b���J�J��FZgp?U??ፍ�4�]Y_�
�ǆL�������BĄ�s�����<����
��g-C��vߦȩu��g�N{(DXr**���[U�*̈��²3O3��G d��rTE%Y��u}������&�
����=�:%N������_잤Y+�����uLMy������,3�.�W�r��q�c�^�b�8��D���
H��TV�{ZKi�j��e<h�@�L�`�!@S���+�϶�ܒ�+�T*e��=�������o�Z} Z�UagD����`��w\�(��^��l�@���Ӊp5�t8��@v��S�^GJӄ$M_�Mn���é$Qw]]� �r�Q`IA��JQBҝ����؅ÿ�/A��XL]+$=�A˿�R"	�Z^ۑ��]�(�^֚�		�f��G�~���:��.���8997��Cd�+**"��IWmrV@
���ȹ�bl>8QN��@Fa��vn�Εݰ��7@��x����g��(���o�b/��><_�W��ŤKX�뷟Ϡ�-�zf����{�B������������Ա��Ŷ����;�?��3�,��0��4�γ�<�}9�Ɩ���5$�3d\�ȶ���?L��W��4d����y�$�YH����✷�#9ŵ���Z����`�[}.O��w�3����
,������n����C��%%-�.���:��x�&�tw��1XYYc�����}����Zvv@�/n%T�qK*I+����3vV5�_��㨔��J�Ji$U�ud��v�"�*u ����7>��	���vMIf�&��N<:�s4H���i�>!!��M�����˵0iit<��g�ф���ǿeX�i����M]�����P�>���@�f�>��1�ŏ=������J�-55��u�6�xr�@�l�(���r�/JM�P?uћ'���8��-���p4�uֳ�#.ݮ�!=0�Vڜ�Z�R��3#DC,@�e���Sy5���uO�%�	B��!�_R#����k�7���˞�I�C�Y#3O�<y	���+kSZL@}B�WSe�B��=_��=���i���0�6ȠOxZRDhvD^�ߟj��
�������������!�K̰�6��5���p16��	�<�e�ϕ�K@��4߿|�:!�8�L�OH��|܂F SWS��탵��|��@��07^�������~��(�	�P.U�I:9�4O�xӽ�����e�RJ7%�Z.����o�G�0�O�Ń�A���	ϳyEw��xZ(����5�������/Xc�ݳ���o��	�+E2��:���E=����LZ���������#�IpC���p�o�.�2�FV6ޔ����o\�MQa =S?3E��x�A@'��NKT?�%D�@�aD�3�1�?�����$�I��xĬRe�$i1�ø��	����O�@?B�5�Wv��yYyƤo��6����XS�fff������t1C�ggᩩ���M�e��sq��
s��
�������sB_��%B�'w.�-�)(��;��*�:��ԫL�(AyT�q�lV�
�b
�#�E7�u �_�]�Ն��f����Ą���	̔ֹ{5��+�!(>�S:��B�cȂ��nE�ax�i��g``:h��Q��ץǆ�dw1��:��py����ʒvpj�7x%H�>��=�� g��L�j
@`J`�}��,������)F6A�]�*�to����� ��ʩ-����	W�[���f�l�%�)�����P��*8��f}��aL��8�;V`f�S�x��]���i�o���TPb�L��p���M�N�~Ka�c�P`ߧ������#�h3i���aojQ�~G�R����k���.OrEjKK���beq1��1 `vD���KLJJI��l����)�`�v�Ɛ�l��$�F�ñB*�C��B�����z����xڸ��p<Zm��T�4}��T�=��h��1�Q�v�׹p�o��^XW�,�xmCCO_��\._6��5�(tO��Y��XcL�?0Xu7�ʶ�A`�^��6���=YI����-�6
��0<�,�x�W�}?��?���7� ����_��r���C�;�桓:<_�O!�����eT�.wo�)bp��|V5^.BB�u.�=�i�F%5��
�7�� ��s�����c 9ME_Z.�ϟF�0�"s=����[�����f��@�3�c��=Y���;��p] ¶W�
2��� �/[���wgS�W�{wϝex�c�?�?��vV&����3���u�����=����~��ޑ���Ԋ�%�����"R_�
3����+�vb|������z��R���Ҕʓ�w�5���[$<��Mg$��y'��5�
\��GK
4�p>^�Vֆ�-��D���Z�c�ϛ����l��oW˫���OA��BRZXG���M�/��.^W>|�f�����k�����r?���m�z����
t ��着"��#�}q-~H=�������8�//�+0��`zU'8jQ�顏���-ő���=��wP?������XB�an����钦0���t�z�E�Cz7���t`E����I����.�+��U�O�Dt��	���*(we���4*!�ᇰ���,����tFy@�!b�}��9�&�?..��a��ϑ�ILF� ���^^Q��A3�3bK;�po���^�&�ԇy!�g�o����~%��
�|i�c��J:E\s0b���E'%E��@��
�_Z��U4��������n�+,�0mN)2j�B�A?���� ��s�R�W�X� ��c�Bt�	q@���3��u~oJ�󔭙�F׮%�ٲ�O��9]������4W7}�PP��֋Ӕ"�� q���()0���k����b��*p9\�vKFS�:>ށ{W ����ONs�.�����}ӹW�Ȍ�MF�6s~`�Ѽs�[	� 0�Z^LV�A_R��J���O3B�x:.��\�x��澹��]p9���l�ٿ�Y��[0+�r�����;�-;`�����,jH-w7b!^���Mkd�FEgţ�Kٮ�����3(W
�������趥l���y�mw��%ϭ��o�rTV�����xփ�Z��0��أ;��G�K(z�ݬ2M�`�猏��Y���.vUP���.Tngy�>J�%�&�q߄��{@m������[]n<M��4�$��R��2���|Nu3X���8F��6���mSe���.X�Y�M_�G��&ߏC�vf�$:��|It�a#{ݠ���o\�����1��t�/^�2&�Z������L��副�����W��{�43���?��MH���+�. ��c��c4!�D����C/��&h9{�w�,,�3&�A�qַ'��o�;'~L|nn��}xQ��7�C�d ��*~	��E���/|*Q��RYvC�[c�����mZ1#{�nt)N�YZ$��g!��L�o�o��K㟷��>x��+L���Z[���?h�~g�X΍@�{�TWK.��W@,
8E�@@��H��OdD��������$�!UUU��A�s�b�������e"��T*{ִGOO���|���(���}�ԙ-�5;���Dvvq�*,,\a�w�"�4��"������V0��	��C-�,8o�Mr��҉RT��
���͵�f{���mddT[�x�iM�J
^���8��}�e�p��f��x����%dc�Tc*
���m[����^2�8w;}��>ܜ���QW9<y�5u��:;�wq��lv�(�Q�;Dطכ�¢�,�􉃝P�v��:��[w�|kv�̎�����3�1�
IۺJ�}��Um�Y�F���n�Λ �|Ԏ�f�_���)gP��3���M��c=<:�[R��L
W[_��?��abi�ӎϵv6gX�����:�����9��Y���+.���`[i�r���k@A%�4æ�jU�{�����0���oD��99���;������n/��sӱaqoK�c��������~�m�����-l��̳9K!$(�wN�$+*)X5i#�-�mA������|;:x��X���t�B"���IF�x���E�N֡�*ӂPPP�;��^p������gߟ}��<�@�Rgk_yn�c��Cw�}�m�z�*�嫅��8F��Kq}9�8�籕�I�4ϓPދV�;���M�`؏�����D�V��+�qX�e��5h�7*�(��s���%3V�{yU����M'��k�j(��d���[�[m˨�]��c�Xf�;�����hl=`�=�Vs}7 L�28��P�)�KV]��ihl^�,�mc��������E�!��B�˳[wkS_�r,��$���h�MLL{i'��_Z�y7<_hD"�˦=�tuQ˙�o`?�
r�(����A�7����B�Ɔ�p�v��y�$>��#���i�G����ZWϤrW����3wǔ��0/�Ӽ'f!�-,�?}!rp�
���+��)�������.h�eD��O!27��0��$~��x���vU�3���A"!ǽao��\Q�9}(����`o^�5����vS�V����:�(����/"DG5��O�(�(Zn�Y��p6���&�,=��+��{�c��dbb��ה���`%'F��E&ܼ)�'T�����#��%�� ��[X���+�~�y�LN^F�p�cC��,���x>�bfc�T�^.p�'6K0�>x�Wo�5w���tx��鰰o��T��I! �_��8�+k�D�M�e��~���$�����;�d�lbt�毤ز�h�T�ٞ��������I ��x&��W���s��}��sw�+�%J�3��>�p��lGEi�==����ƒ�d�\7n*:�9�����ͤ��e�)�>���R�Ң����dĞ�IHH.��E�S�ړW���~Hf�� 2!�!���!�fg;���{
����h8�@����d,�8���W��#�yH8��8���ISWڢ���;�h�Գ2KࢪI�Q�H:,־1����F���b���\�y�� |\����j��|��O�]�4�`�A&+:c���4^�Am�s�8�z.�g�s����ag��n 4؄C*'D�"�5�#�F�I^O�HZ��p��y��>�n����ouZz�U;@ >����1���-����FF=����,xxx�\�􌌌����#��.���&�D�5�6S,���o�*ô~����������w���o�����ihh\nvAĥ�����������IF�? ����4�Xd���y�3�V�ͭ��ƪ������UX�6�i7�j��hJ���d�̦,u����url~2�HKG3tu�O<8$�A����s&F=�����ߟ��H?y�*�Ho��0C\~Ar�Q�V_�*�Εt��lLfcDǋ������B���J�Bbźmk��zF���׊��B�=KK��b6����������J�o��W�_;����z�67��.��d��3ܯa�3x7BO���j*kh�y{��d����a�����u� Ԅ qB����9B=��F�=���)A?�����	��!���|�e\:=��YV��5��t=�G��F� ���`�?��O�I�j�&��Z��Q��廘���Q�lҢ�|*����k�Hi�7T�L�f �A p�}��^�v ���[�Y����C�uGƸ3�ce�{Vd�k뚛�IN  D;ώ�jj}�e�-� �#����t��(Dt$���FFF�oh�=8t���Nx�\�2Z��}e�G���s������^�{~�l��-��ʗ�$1Ϭ�۶���!\W������vY-�?�יa��i���*��uB�QɃ��Uo�UԮ?4��Jww��!��J#� )�"-)�]��J�4Hw�t�k��|真�с��}��Z{��rE���� ��:��,���2��Bxx�8�{����7+��ۻ������P�N�v���%��ߖ-���UTT��k�2��9����G@�xnfFs�7�u!/'����֪���N����&�S��Z-����EJ]���� ��aT*�9��\m�G�3tVA$��۽b��<���d�
r�_��K��q��A����N���������fo��2J鲼��Cv6%+�oB.�DWᡈbW!�܂��T�aRV�}P�B8CCCh}���rv��`TDʖ�>���ш�{Ӕ�梔ݽ|��.�-����w�gz޿{r���և�OGG�"���Ӧ�=�=Q�	��'�/��Şijj����{�cS����$�∓�{p�V���j��~zˍJ	!��;��������ã�Ԭ,���K��<�rѐj�zSSS:Fƒ�0��X�f�sY>xg������l����2T������j��7�x�2z�%��'���]�ӳ����-��Q�.�1�c	+3��%�F�9fWw�n���s���  ����i8l~�;�򷹠 �����w�[�'R�r�e�ź�1?9��r�1Rz�$i-�-����-��j����[|�03��`�%�2�Z���,��#yg�<�4
pZ�C᧓�
+B� ISϿ5mrE}b����B	�/��m�>�N�\&�:�I��S�������� ^%����H�>�a���8ñ��	��77F�v���Zk����ؤ�&�>ߧ�Ll��h����/��n�РSf�o۔Խ�2S�tW�i�>�Z�l׾~(�-��폺��(|-��O�ի7W�+,Ƃ��t�D ����l(�g�=�$N�R\?��&� Ѝ������p���	�A�!�<��Mӹ�F�pz���&3xKؼ�ㄲ�)#����hn�S��ÿ��� Ť��\�A��򺍏�.��L�Q�;w�����!G�z⻆�˗�B�jG�t%�����_��Ǩ$%y����<������>sI<�+887������BƁ߻UG�)'��a՞�!d(5I<�~owuQ���6��8��Ă�����767i��H�����^����4�q	��|)��{�������f��ob��r�3jvXQ�<�G���s�+�ns��,�@a�p�]���RE��m�(�~A�?��'�am�yrh�.�P�1����[}!���cu�����Z�D���^�F����<���I�����~�1�Ϫoz��J�k*	��*k\����2Ѝr|&k��:b���FGO���K:�vzz�|��=�f�N����;��_��f�?m{NדUY9���)>_֖v�^��ż�,2,�e>3S���{�g�G�N֢��we߃�c���i��g�Wx�n�[1�0�+LQ�G�v�eddBƅK�&�Ǜ[C���D,<��dx	�;C�yR�d��;��y�!��Y�*]���B@�_�.�@�����R��%vm�	^��_�
+P��}�h~��S��lH����p�(��˿�N�S��ETP\\�B2�4~u?��pF�7��>����`��Ħ~�%��7�$n�y�nv
���D�W�
Z=��N�*}����<=���[0��{�V �efnni�q���:�t�D|��A43��]_�s�LB)�`�l����o�yY�ϟ?/���ߓ��q9/?' "i�i�^e@x[�fJ���#�i�ZL��MW��|;�h�<�<�H�����4]��$�!{�~�����G��\EZk�>kG�kĊ���@�NI=s �P7�on������A�R�	�wx�����n�����ɒ_ �f?�L�����^Y�vl���g�QS5����_���5��Y.�R6>��M�=wo蛯PA�+\����Y|LG����x��䤏������H�Цs��Х�Y�˻7�L���b�#�U�\'5�|�:_�|�+q$>�ҳ�`bb�l�F�pKm��stC�.�������tTj�*}��d� �������Õ�ݞ飦�����)���s������>�憆�Q��4�ɞ�J��"����Q��¡r�/�-2䰉�
�-�Ӷ_8�rħz)��S�#��z�
:s������Ĝ7�3�oМ�N~y�|���.��ᱧ������o@\12���657Ӳ�c200�3&)ᒒF�p�>��:4�'EF��q̒�I�h���S,��k�(�G�~��,L���z�y{L��w�z�{5���`%��ʲ��lm�MW�X#�rSӥ��O����6�Vo�F�Wo�xj�+]��3��\��(D�Q544X�fj�����C���6>��6'�ۋ��6���2(<<<*4��)���5K?�ٛ��?u��_M�<T�����|��	��� ��E��bb�����_�o��;3��O= ࢢ�w�6��"L\���]R���(E�*�t!��_̳���sv����˻�fj�H\ɿ�����ӺK����IC�76�YX0�7�8��BV���|C|vv�s����V����o��d��&�_y�iLL��z<#"
��ӺW��Obu�؟��S����2��
!�˯��y����'�l�R�7���p��H/ԕ�b��������M�|}��{�!"�����N" ������#��ouy�C�d��<0�x+���	jjj����m��F�j��)�g*���sbk�3u���.����pBζF�&&�7�{�����I�q5q��v�ξ��ccc���զ��ag����++g���錐�4�����yoXz�K�?W��� �UI-�eQO1-G9
�E�̓����d�����;;;+@A�;l�0��EtMM��b��_�d�)ڼO����Gѽ��o����|���$W�m�}R��F�?1��(������}��w�(Mʋ����g`�f6T\L�?:�ܸ���Z[�.�F4�����Wk��;Em7�Gm]�G�K�|󱂰�� ؉h:��3�X�0��">%&"��TQVT��`�c7�������WL��r��@Y�J������w�7��ɩ�5��_	�[cc#���� :���8�t"��|o����[�ӛ3A�EG_y��Ё2���0&������H7;Q���������JØ88����[�.�����E�n6+����nʷ���@��ܰ+).�zӉ�WX�EF���O�\�*���/W
ar�ru��	���9M�Ǻ�/.<�S��������^wV[T�Y��***~���qp(��y�N�'�M����h�`R���++��|	����a��o��C}���Z����z�6�ݥ��Jy*b�9=� �gm-�`��چTcU7��p�oZ"t_s����G��A��S�oWBb�m�*����9_�Z
�?�*2$�y��n�>���?��:\lEG@@�&�Wڰ{JA�p�M!���9"��{C�9%��@��Z$A6Π4�y��B^���*	���20�o�����X�o5�E�2��Z*>�� ymT�!����8:r���sA��
BT�TA�g ?xq�3���ӪYY\��((�T��t<�& �� �t�V7j�k���Xh{4WW"�W�PnҊ&((���T�W����@53,C�-���QLi_>�����w�F�#�gg��l�����N���T}�1㦡�e�jT���˰�u6}�v8aԗ�&�YEY��s���ލ�ӧ�b  ������?1� ��\�ڂ�y`J���!��ai��>���fJk}1����-�'s!j�����Փg��&���Gvî������=C�-l�E��9�cE�-V�����Xu� ]�-���ܮ��m��>[��	�_U:2?��>W$Zp뛸��t4��ߥ�&f^bW�[���J��=��N�����|I)�c��KB���3G�Yd���n�!zz£X1g/e����X���F��/v�Ў	:�a��G"�?�F����V��溁�;]�MNN^t[\Rb�ׯ_���,b&�H��[�_���9�T�6GB
�	\�6�}U�ި)C���n�i�d� .�b�"C�*5���#�^B.�(X!�U&�c����[hrC����?���|��om���)��fN�`RY}
�-��,---ˇ�X�ߔ񓚧�Zc������Baa�]}�O��s0a{�YW�i�6���"��T���������kt^	�����_���r�MM����]Q�'�t)/c,Ӈ����'��iG�v|y�wu�v=����7�?{y�r��������驩��|\B�P�,�	�)��\����Z�7��O����hxY�r� ��lm���˧m�{y��o�c-#�&�1�&j6���/�U3�jiuU���v⼕�H�qM�I�E�}�h,�c�����E�cַ����[����[��ÿ�|���L�� X��������l� }�H�9'F�o�枪0�t�dW����}���A,����%-_��j�.�������y�{��XuK?5�g��C`���}G�\AT��r��q9ݩ-�'��'��g�d���x�ܣ����bYf�0��X���U�0�k�J�|��	�荝�Y�M�9/>�=���ϲw�C��gKs{���֖�m�|zzJw����O���,��_�S�Yo�����#�b+kb�i����m�����596�F���~�c���ie��e��:��U���>����NвEZ��@�h�������#��*�M��3y���@o8j�S.�?�z��ip�b�JXjOOO��n��Z5u�6#4J��� �HH.�,����1aW[U����^KӈUz:ˎ�K�o���[�눜���K�\���M���D���$���,�� ShO(�a���*�e5H�և��Jp���y	3��(��ƣ�\��9ƀ6�P���[��^'�W��â��;�uJ,L*���������o�o''�a����D��ח�[X[����FEE�T�]'�u9l����t`$0�-�ru|� %QaAMM{qq������(�����;�d���bZ�Ɓa���U������a7�d[��%��yV���w�Bڣ����$���@�A,�a����DБ�l���<�������mk� 6�;̸�s%�2��;�)��.GN>>�d� �^��c��;����ں���b֦M���p ���H�p�sDa��J��)#0�VG׻CXNnn���~��H�]Ft4������K���mO理ҧRXQ4��]�Q����]I%����F���or�i��,9��$}N�~oo��X.���`N~>R�{Sc^����I�DJ[��A�#����D�!qhh��A M���'�z����L|��"��fll����$nJ��@��W�Z�ugw7$���2(9����?>33���-$<�VX8��	5����ǜ*��)�r�,�@,�Sb�7��,,,۳u�aXա��ˍ�?��cx����Y?��������Y9<��H�y���$#3s�����S�x�x�������w����X^^^�9Ex��E#cc�i=�����׏m�d.0�>z?Q$�x�,����LO����O�t.�)�&�hn�I���cX�@���n��y`j�7Z�(.����G֪dK<uqq�q0�~_SS���� ���/)�0�M�������k��\-��]�G���uXl!}��i��9�$�ۋ��'�Z��sRs�U�r�&x��m���[��CmZ�X������W5�qC�����tY�~Y���Y���a:���^~z�&��T��$<�"������q좦F͞��������g(曛�3��/����$��S�����y��ܾ�޷�ݤ����|�V���y���T����T.8�����������>���'�\Ù��^�4�v���]"a�<���K,HJ$��I����H\��lOǳbw��.	A��bM3���͛���9^G����ӣ��3Pqq�����!rQt��H�> K.�&w�ֽ=�mem���Z�O���nx(6E�h��QJ�H&�k������܋�nqJv�j�*�=���/4�'''�nhE�m���t���<����WaBh�������|�9y<]]]&�yЩ�_�Q��Љ�:zc�e��^��M�yƆ� ��P�H��@!��ɻ%0̀$�ȈZ���l�n{,j|�w�o��J��^�����CH�ooo�t����ᅎH�|��kd�:�kփ��������U���'F&���2A`W:���	��_b��Q������5��fre�[ޝ+m6��n(��7`������/����|&F�5��"����Z�i@��.���R�,�J)� ��r
������`���m�eHh��_=cc���o:��j�4�/4MXEs��Et_����5��k5EJrA����[ffvve�+�5�l�㬧g����_���жQ�wu}�մ=@AE%�.��cd�P-;�&Φ7��֘��N��c�����5M���:�/����ON�1��穨�2 W�ytQ�fS:L,,9����0d�8��-�?*k�su��n��/> �U`ˣ^�d�F1���iQ��*s�4@꣓I�ko�¨����f�M��;�H�p��G¡�34�3N���ܯc�h�T��%�\��T�[ۈ�=Z�C�-K33x�Q⾺��t/UTN �Њ�Q�V�{򩿛�Cx8JFF���۴��f��F�J���o�&�'�����G�}�&���Qӄ\O}��)����EVBь��Cp�o�b��� +3l(V��F��rDW,����k�h������l�3���л�G����?�@)�Z;%���5�{㶗����P*���qHHy�J� ]�7Dm?�W8�-��4�k�߱���1dedr����Ḍ�-�f\�Udh"���7�v�$�H7�|K�(��obr'(���~�e�w��Gj�6��i��p��c�l����/`��/���l��9���>�)xl-��K�*naN����j��p-��z��m4iii+ Q�9P�������{�f������ߙ,��:A%��U�7{�-�W�K]��MsDSkX�J��cC*�w�cx_7q��F��N�i_;��ȇ@m�rU��Dw���c��U[˲t�ʦ�%Z�X�e��c��M��n�o���C�0Un��G�z��܏#��$�9�)|�x:,��F�=�����yr�~���hii����V�������s��0���7�$����C���1T���s�Ѐ&D%��FQ/ʻ�N�YɧUU�x�jJ���ג���C�בI�Q�۷��s��%�@*D�����ڌRMTp�xR���-��?���¨�O�aɩ�>`�뜛��3p>��Z����&//5��ׯ�T��h���%� �qm�*7n6�A�k�}���h`�ƃ	.Y$`��:;�'Op_}�WQ����"qgz�l��s�I��jeo/ja�(C\YY���U��ρ��P���Y ��8)Ɲ�7��^8��X�i%�g?����#.-����^Ǜ� W�W������hŒ��6�]W���no?�xD�7�Nmp�Q�V��YA.t�gfF����@���)��p���c���b��rq����p�y�	dwtt���~�gB�
�pXG����^���V#�W�^�@1����B���[*��Í"�'FR�i���u0��F�鴘�|�S1�i�p�;ˌ�۵$\TDY�::zәY������:��4��{���xp��Y��a�HY�����>>��xO����d����0�����]G%ی�½�}�H�}�N���ȩ9�.���n~}���q\��Y]᪚-�%�V�����í��d���즻�U��_��<�w���3=;rي�G��z�(�������5�lcB Ļ[}O@��	��gSt�v�Ň���H�´��q����]�Z\111�8N^^�������l���
E��r����^�c`t��+���ъ���������wxZJZ�����l��Į��lD���|�����Y �R��$�?��5��F0�l��� @E�䬬gDFe��"�y��6�����#���䷵�3��wH�(��"� I(��Ԍ���U�{�_�
��v��S�Ș��w��,>F*vv1V@��~y�mI��J�;t=�Pf���"-4R5�k�|c�?;�7�6��q&"�CP��"��G��]9B���O�R9_u������}��F �e{hJ�bN^��w���,�j�����SXr�p���:���ܐ���ŅĄ����z֢��Y������������-��rsq((J+���m��"�B��r��_�R0LZY���`�(�e?���$����m��� ����ŝ������2B�N<����Ӎ�ɫ;YL���'�~KH@�z����&�зc�����t�����$�|�5�DG: ���o��7R��T�����2̚ՙ��-F�(#���d)X��Eު�MNB\�I
5u�]���x5�R��F8��2oew���=�OI��c���~�E�ýSF�����pU��6T�,Y��xV��	rt{�r�f�(���C	祥��7RLu��|�E�5KMV�E���:���|��� �CA��[l�Rj=%��M
2��ܥs/��T^��-�������:�č"~�n_��ɤ{mar}��59��O(X���9�ZV�Օwh�+���"j�d7K�B������M}��G�h|}O�9hʍ�)�C�S��ʚ����u�I|�s��o߲D��H�ZZY���)�1�;����*��`���p��v�-,,�n�X����_7=�d�zq<ܝ����� �T�o�yI�3;^�I����#�䧵�k�m�ޜ���iji�5���XRj�#<���d�'����<q&����_n����5�����GEE�<r�iph��|WG�� ���¢c|og��UN��� �]�NR������	}N����tޠ����vUD��,����d�Ί�_�]HXߪ�M$a�K���e�|����J��(\����쌐� ~a����x��#?��NIm�V.:�ѩ:���gWW)ĩ
�8�����^��xO(�J�[�$�����\6n��{ugK�C�®m߭�zR6�.7n���(/(����L��fL��K��444����:#BCC��ܺ����p�_]5���r�#���Md�:;Xj7�6ף�������q8ߛ���2@J���(����=���l�-q��]!��^��v�3d��ow�999�����~�sP��~����
�HE�*m�0��^����ih^����^L�u���\�������\fF�:G=B>��(	B[A��HB�U[���ļ��m�j5�-(( �������iQ ��!7o��˚*�Ü�$�,f���]����a�SRQe%	D�n'p.d�l�1I{�������y3=Ħ���%P׮gf~j�;7��
x���`�,�7"��ۍ�u4�(Y���!�mWR�k���V:C�=<z��
+]���S��y��5%#a���T������B�Y�|�rw��:vqq����<��ѥFy�k*RdP�=���%�&֣{��qyf���͡=�#666�zG[e�� &�8�.^�eU��@�JR~>���q"���ȥ�%���1�V>�c���4��(�|Byi�B�Ğ:�Ij��6C�v��=�_Ҍ�#o��r���48-���)���g���OEA��}GSu�Eh�::���"R�� ���P�6�x�XX�fS���Q�Ej0����pqq߃X�h���vc�=�+�uE�ё�j0�}Nh�(���lll��D�3�3N�@�|B�"1WP�.��\��6:5��9�.Es�gK.�t�c��lx0`�;�
J�;�C�[_��I�i���&�o\�Ezw���r��+���kk��,�m?�_GZ�nK�^�}��(���G6�hԖ,�|�:=6�@�����j����������zj..u꽔$f��|ݭ��hz��0c�Y�ۻo������-�*"b0:��_dgg��x�K�K&���R����͍vy8׳�G��M"*�5�q�OiI%���}@s[���.��q���H�.�.�s�]7�}}J���Gh��o���`ߴi`�^�/�C�I�K{���e����siM�+�d�A��ZX��w���fѷ����](%����^\LCK����C�A�ﱫ���q@�
��L�4Q��e���xaT��蠌�x-ZV��(���`}e%�\�+���ly))x ᒵ@�c�Q\����������������𵴴���!PNfӘ��lim�)�0�g�gt����^E;�����j�XD�����#4�" 1��$14��O;Se�y�΢���QO#�ހJWK�^ݗ�oT�X��D�7��#SBTDx�(--#����\쵭�vi�C��MB*�ǧ�n��Y'D��~�
ס���C�8���6�T`D�+_�]-�����`5k�SOFK�0�-��Q�n[XZ� ț;;�KKK�K'���-,,�CI�������/����NelM��n�hkk��ۗ��>99y��S�نNĶ�^�}��vKOG��������ɒ��		���$�����N0�����11��<k����600p�s 0&��<^��W�|~}���.��RVv��ﭭ��kdT�������t�����z�g쯪C�on�w�ր��x�E�]�v�����Q{�I3@���g��6�9#�ܾ��٠4��=]]W�II���K	s�;���o�}ss���[�2��&7�z�>����|5`Z���ݚ��� ~�@��,hk�1��������ZI�7j��'P���2��j����T�%2�[���|?eg��tOLLx�S�`wU���f���� ��c�oD�܈Y�T�x�o��Әg��}2H^hh�4,,�g��U�(���I�Ҡ�^�yC��Śd��4jMl~��q�����h�����~�������З$�6�K�(U:n�x��������e��2��׊��z���)��
&$$�}P؃��&��y6�-�n^^�#Y�Zsg#$��w�_��H.�vRv<V��)`�A[~r��%W��>��J�'���@��� 0B��Ƿ~�r���~�Q�������`U�o#5B�<��C�T�L��V����'[6JJ�x�&���P�$g��ا�������i_�(%.03Y�cccWm�./��}��{%ݩme0;)�~�����׷�33�n}O�ԭ~���� ߟZP`���ވ�?�C�M��%��9M���JXl�&  �\�p~��W�������ן�k���[f�$��6��j��	*3i����{��8�V�\���u�-���z�p~�G����Tq��2���s�t;���9-f456VFs�*�gr�vvv��|����G����M�X���u=�jr^	�O�q�Ыx����}��Ǫa��\�������ш����t�5���}�b����ʠ��?�����)���V]����ٍP�+g↌ፁ�y����Fl~�N�~����ݐ���	�O�hIX����T������5/�}||�W{�{zB��/�*J�̵���z�����(J��kA/�n�'�.;�6�u^�=}��*�+���P�����Z%a�$E%%3		���ٴW��z��-�� -Z�Z��R�o�[X8MXXX��$��[1�S��&N66���^����3(/�K=ݟOa���{�z�:�Z��O���]��`[��ܬ�����)⾝S��>��5X��y1��?qү2�M�S��gi�<�k�������}����{�k����e��PJ냾 ��U=I� v�K��݉<@\W��W�����Ɛ�=��"_��#�#.-��G�]��O���f�#��Tކ	�<,yo���ܞ�Q�RRR�Ϫ췰��:��~�G��u��U��q��xee��0LsPFV�ز��Ǥl���g���4�,�i�uNN&��_C�OF+$��h`�E[���f+���r)��%��A�!�����}���第a��������*�N�2��.,x�~_V�0\;^�ʘn�mwbM�p�����_�N���`��l�8�Bff�p
22˽��L��"��-J ���oKkEW%	���(%���_�O/Y�}��m�q��=ȫ���}���^ȦUVr	8.4�:�N�S��fl{���l��8��y˨����hR�m3f�->W;����j۞�����#i��Ƞ|� h'��M���.>���m���|fvbsss>�9��@ߍ�ʢ�v�͑!##+����������Cg���L܊����{�`���Mz�5T�s�*Lh h��?�_
ŬF�b[}���[ߝW>��xE�f2���i*�����Я_��(0`�;���ñ)崵��� *@.��PU����_��w�4yL��|�
���P���L@@ �}����3��H��#_��N��ZZ[��c�t�S�M����yB��t,�\`y+;����&>�A|�$�/;B��K���ӯ�G�ļW�bF�� �'5==�{+��F�A]0�*@�2�6R	m~QH����l٤yO�Rͭ�m_D �|}�A���i�>S�@���m+�`�E��X�����b�Y]K�t�Y\ܘ���Z�����W��
5���		9y��d̜���}e��|����YYY��q�_��ş�N"�jt�<6�ܱ�1lK4D�1�����o�b�������"Jy����UK��<��遶�AYgdd,C�c�g����������7X�����|���-F�<׏����\||!�4��
&&�B{ e@@ ���BSMg��x�]c7����rTs��%�B�?������\�����]Cy�|t��_�W ����c �.��ɐ��s[rrr�Ąv�y
P���Ԃ�zyq�Ż�ٶ����+�tw#���j��1P2�ЉFp�~�Z�f�3�
��'� ���f�Я�Բ�(�3���ssqy#""��N�ԁ�I�}����Gmg �� P�Jy�lv�,��i���uX��/��a�R'_�}����OMI!��>ͯ����\��P���z#"$t�pe�H9G&贸�rA��H���M�I@�$��FzK����3<�L���<vS�+��n����Έ���~[�131]=����\Y�	z(�Ց>��lSesyY=��/�kT�#���bsF�hb�pqmg�������̧��~/ɒ���B�c�:�����HJf%����x�8$0�W�V�����މ�OP��5�ֲs����!ڱww~�dn[á��������NnFDD^��uC���jG�1F*;88��1���:0<�FYM(.7��_o�s.O�&pY���XM��`�w�E����'�����>{6��o&�qo�좀�[�l��5	L6����Z۹����C'aG2t?I�_����<�VVV.կ�wqq�+��fai�fk8j@�1�����:��Lг
2ss��8��Nk�^�ќ>���*�<;Γ}h��s_�M���,t�T!`����=Cf�ӋUGG� �8�/#���D
j��q��)�
f��nZ^[C���������G��!j������ߒ�R�( �h�Y�0O h���)��2�6�'^^��{��@�%�<׃�]��$��/�d�$�)��_:��N�z{{��,�!����Nm��o���K�UT|�aچ����/��+�a�^��@Z\\L9G�����mU�������1�p���s:���GGq�����4@�:;sm�yK)l�ac�{{A����[F��ODP��k����@���IPc�����2�>�R�<<���.��fkikӝ ����f��넛�r
G������:##
�����ƭ�?n�<��)��R��cSJ������x��3�'��lu�����\V=�B��N3cK��aϳ;ph�T`Yˁ��i]�U�K˔���I˩�f��b�)�>{?.j(Ps�\g1��%6��F����Ύ�OKR]��+ �5yyt�4}cd@��к{x�UTT�d�K�a���/�^�'��Hte�և5.���$��g�ߓ�5ǿp��:0��p@v��o�";!����/[@)�L�2d��_���{h����~����p��7|�b>�ݾ�ǘ���5��>��L��8`0�ea�4 �V;�#@�����@s8�����]zn.t\����f<�	4=RSS��Z�׉khh��H�g�$R��φh�0 X�e��������?���Iq�$�ccc�E���'��o#�! ,b|�7�-p� �P@a$�HPO��
�v �(�)�����
��wX充��a�x,:���2��,�\�����lciYY�높X�]�Eȕ�����������Ԏ�a,,��^i�r,A?aS'���qh�:Kp0q��Y�G1 mU{�$\0999!g��2C�=�;Uհ�8��ا�@nB�?���
���$֠q�G�ӧO����gp ���΃&�tӪ�D��q�kmiQo���w���ܑ�n�J��k�h_�������tC9^@\\�}g\���o����Ĥ�猁�����·ͤ%5�(ďNL,�f�cX22��A-9~ls�ጕZl
!u[7�B��]����&�nxRo�GG��L�(����PvuuEEK��h�E�J�ԃ�#�tNL@�u���/v�oD�	�8�2Q��_����	C����&��pv �ӧ�I�ʤ�]�PGFf�f���r�Dr�mD�[��\ R��D�&l�/A���3�o�Y���̌���:��F�m����˗��m�[A�sRI	���5I�l�ޙ�����>q��a1H��|zK��n�s�g7��;��7K��a�===3$���^3���]����X���>� �@Pp��Dl�ղ,~���q��cd4�L�]7Hgo��V�.;\%\2*5� �s`�Y�Ag~����8��k���ҖcDw__`FPQSUc��'��z�s�o/2�C?|���{$[������/	�.+i0Vt Xf���y�
�.0v�
��$}$� �t�)pqqi��z{�}Kcb0��F-wc�A��S�&|VjԤ��������ɣ��O��2�M�7�����.�)&de�5#�����hjN+pb�@;�M���eEJJ�ᦥ���pi�?��/��VPX�w�V�� υ�7��&
GS� ;�B|~׺<i���M(�l@�e@>���}�r_�X���2�C66��4�.)I	�ru�D��b�TJJ��߃W!%�잆��� 8:���`0]]���j����C�!�x�L�P ������۝Z�!�j�S*^���N�V_��!���&3��_����N��d-)9�9�\�5V1װ��7]�`����3�%�E&-��϶F��hiqP+y������8^k�'&&�]�ߠ�.� ��������1c$�x��Cf�}@��*�Q�e�8MۺA�T�Z�v�!^8� `���\��)G������;������sHH���uR�<�3^�K؎��<��.3�sb�$�~�A%Q ��i�?��w�V >�CU�I�w��g���ꅪOmll���"����`@��{���ߊ���}s�����TS{�aff����9�guzqA�܈M.�a``�}y���C�Ǐ��((z��h��~����,<��ciħɟop���E �J9�����h��k��Y7�����ÿ��� �-�q �������AOD3�`�8��ê'EE�����k��߀�:fH	��+�nl����K9�.w�AOMH}U?F� �	

��;���xy�CS��(���=�Fs����%((|��.��@Xy9ǿ�sȻ`b�`���L������F���T�;��ʿT�Z��Ϥ� ��ёp$�Z��k-l����İ�c`` �i���xf��մ���N�f�PmR�Vן?	gm>@���%��LDD�Kz�W��`/	RFDFֿM����ҹI����p	��F̭��?��aJ�g�V__/�I"��}�����gK�O�����m��F>�B�6�ם{NVC̵�����F�$T�M�e�e�+If�7б�_���o x�8@9��jg!X�;	�	���1�q�K9X��n?��Z��W��&�[���(y�?W���ju�L�q{�f��N��H�e5dƭ��`^r>���w����1[��O�S��l�
~*�]��6���q�?K{!�\�rsǋP��t�O4tta�6��X�����i"$�%���%L�H�Mz ���Ȉ�i�����Z���=����cm�����NRp���pQqqķ}��kS $�w���ں�V
y=�����86~�$^U����+��������%@x��w�3>(��픋!�]��S�*��E�dm�R��Z��� �4����x��\�Y��ϟ��*�����0:Lb��=0��Z������3EͲ�JK��m�h"���	l�ϙU��A"��w���G�!�j���v��l#�0.�%ػ�i���^��k<�J�� ��I�l����&-����N�̕��/�m;�z��@�"�2<����{ p,,,�AS���K+)�����E�����;�����Z鬉���d��Fd�0�m��7�T	�
�_��Y}Abdd4���)�k�/.>11���.�x ����7��g�������!Gʡ�!�z[  'W'�Ѳy����Wa����l*`(H�̄^���Ә�
X�ׯԀy��,2:6v�淪%��;�d�=_��� '��p� H�O�AA'��ٻ�϶\�e��h��I�H���F�RE�D�p�ϋ+*� �z�'���*�fn�*j���Ww�P��G�H�e肂��qq��o����IHHlH8�����V��2��z�J7�.�\�8X�����pn���|�������^#���P��$���_h��������Z��3�����v%d��T�Ԭ���UP�A_&���T��hKOp���Ya��á���������:������ϼ�g�C�~~bK�8�e����n]���f8��FRB��<?''	���nS G.4�������1΍'t��|o�5N^�!1>�����������'���ؠ�m(������o��A&�����ŀb����r��j��}�f3|%�2Uʖ�G<������_W���O!�@�)�*ä��B����	E�"�E-�o0 ԀH�	��@)��[+���VЊ@�P�*Kz�t|?ޯ��sϽ��Μs�2G���J�0E��z���^�����˹��7]��6@z�E���f9;;?j�� &G��תa����S����)k+�rB�������M����*L ���[1���&���O��bg������J�Rٔ��-��D��I����d��K�^��S�X�.y�m�=W�n�x(�nP�]G��c���l��ޅ�9JA{CC�E�BI���qrbe)'6Rz�n��VT�(?�;�3�Ɛ��Aa(�/��:?Y����a*��ɣ��11�����;;7g����r����+��夙�9+�h��>)�� ��j{�?-m?�Pi�	��Ok#ޛ_TT�t���Zk�1�
3�G�gffy"�oY��d���8�NL�'��'�t2���U���"ȣ����ܟ���;F$ABBBq�DBFD����+�Q�R�٣�4@���79:�C�!!H| s19���d��+��;����$��7����SL���!V!▪('�v�O�ʫ�"����􌌌���Ђ�@t���՝C�ҲX�]��f��YbRR�L�/�a���{]\"��v�%#�-���Vj�g�%9���k��3'ڡ��zSQG.���);P�~���-��H�5�[�3��5d��{��gݟL-��|)	XZ"�o����6�+U��a0�Rd"MX�T�]<�R�+��K���̒�9����m�9~3�e;ɞ�P�ȴ#��5練�;<	결d���K�������ō1�61�}!J�U�=E����$5{:��Y��$'M�G{��4YB[|x��yG)š,<.�*:��\O��ZO�g~�m��?kku����$'�I�d�w ���O�\�˃�YG�mrH5���ax��Os���w�B(F�9hb<*4g�	�'�b�d5'�m���Z<�QM��Ù͕v�����
u�h����&^T0�B�֛�P�t�ӽᥪxyu�6M��p&���Ué_�%�Z���,�p(�صM���zQ���ź jIw�u96���n����h��m}��"�)Be�ـ͵0]� 0aaUu!�4��vmi�cȥT^G�� i��G�RL6.{��*�\l��WTjq���3ُ� }>��9_��PK   F�X ��ɲ,  �,  /   images/c14208cd-713a-4fdc-8661-253b2f19f73c.png�,RӉPNG

   IHDR   d   A   '��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ,:IDATx��}xT���;�I龜��z�EDDA�(*��RT�`�bGAD� J�"E)" %�B	)���}�L�����dD���=��-�Ü9���{���^{G�[�F�	���+���h)�/���v�J�"9.���r��2�f?�A&�ޒπ��h׮���PZZ���x�8qEEE�?��ԩ3"""������r9s&�ӹsg;	.��#��E}��Jggg� z��>ݳgOL�4666��r	E�y��z�g�n�����]X�`�7���3\����U�3&<�{������HA��M�0t�P����gϞ��Ѯ:��Ɋ�����J!Ɨ�����Sp�=�`�/?�Ѷ��t�CE��c���b��4 ?��&N|���V;ڻwou��ٳ�8	o"��8��������z�^}��������$X����,4 ���77'��{+���}a`,\�5��r�˺o��� �F�pqҢ�$G�Fa�=^x�t���}��h!F�����m�!�`�t���c�B�>������ݽ9PQi��{��1�F���G�����?���E����1������������7�`����׿�u��������x�o��ʰr�JG��_DZZ���q�w"55U!?&&���4hZ�n�]�v�C�عs�z_�_�^�[���]�}z�¯;�!/��|�Ĉ�pE9�ЯgGie����qqq	���n��ql\� �}�&O������r��l�A�6�����9r~\6��F�WJJ�/d���$�[��):��ö��=s.Q�Y�‹s�Z��f͂����WWW�t�����۷���|�%�<'A222�p��Uċ=c[-[�ĪU�Dm܋�b����>}��"!>1�h{{[��]AaQ��޳�>���\!�Ytl�\�k�֊���ztmq��$$\����z�#5���m�v����~����oJ��	��V	"7��G�q�ƾ�;бMc�49ez�}�:�7WG\�����v..2"hDl\��V-C9px=�RF�\޴iSš�Nd������ӷ$���|�r<����:�ܣG���K�C�iԨ�RqTI�	x��5 ..�o$������GO�	��*����5�w�lFb����C~>�j_T�U�j�Z����VZV>�Qc��K��~�wm��ό���^m#}�+��e� }�Z�pZ+��̓�P�����������pJ^}k)�|e$��p�t�����V-����z�j�1(,,$����l� ???4o�W�\��>�JjѢ��ڄ�"�gΜAdd��v"xԨQJZH��#G�߰�ѣG�ȑ#�(�cǎ�ѣGQRR�r:�R�k;v��]����|���+*^_�9�*\������������3J5����O��]�8����ё���fi���#W	�-u��AH����A�P�>�R];E��%��F���o[7a�˯+���'R�$ڏ�3g���?W�(%%�V����TG<}���씭ؿ�����:u�lԷl٢>�����P׾��[�a��!<<�WSO�^��g�����#�k�|�O�=dV��Aj���NWVV������,�Y� ���J!�VkCV.�.���v=�ƃ������8�3��"�EJz�\I�pW�d޼yJ�����g�ƃ>��u}HH�B�5��J��S����;7���nd���2�	���o�N����Y31L�&8�hM
��2�N����P�&�h�l/�������JJ���������i�-�3�����/^����%����O>����F�j�*��ƌ8w��}twM��@��5�������~��0W��.���&8��q�g�z�����\X��JmTi*�q.)��〼��:�C�%�%��rT�@8���iK�\���ydf��S��;z�Q����~�V����n}ðf�FL�6UyT;v��w܁u��)o$))I���(A�p�}�������A"�S:~��2�?���Ct����gQ���|����������|�������G}{����7����!�,�X�s?z׳����J�ۜ]PRZ6��To��.=��`50ܾ}�� �p1v'Z���W4���sVnn!|=�3�O��*;���旔����Y�WW#QD>=,~RJ(!�.]�C���ݻ�s�����UH���QAc�����%���>�O�G�1BCC���e˖Y�?	d���"Ti�D���(ӗ�?7�4�RY?a����i�����'�U�^ؽ���J�5kV㡇FL��؈��{���W�K���'	�[��p����$�����1��ix�w7I��ѣ���O?��?���7�z"�6�b��.�'33S�5zc�N{s��u R���H:�J��w>��Zm/�mS��1���V��7o.>��#��~6�������n�h�EҿMr;G�ZTR�����k�s��k���"��3���*A(N����D؋�q����%Bb����`ޖCH���9�>�FLį�nU�Ɖ'⧟V"�R
rR����c;ѵ�"%��z<tqyٖ���+��$X�V,�i�H>gy����_o�9�M�����|elK������Ǘ�|U����_��S���W^��e`\�`t�c/��U�к���������M��G�\�e�9cԣ�Ec�`vTn� r�ώ�'�~���l�8�W^_(����4TA_�E`P�;F�\���I�&)Og@�6�� �W� ��q�=s�xj�U/��E�&b,]��%:��~~�
h�קâ�K�������L|�l'�<;�g����{� $��VU���������Ǆ	Sq��D����:��F_.���m;@7��SM�i�z��;u���Ga���bd���&��ؠ\���a��O#=?���]�A��u����x��nA���1�*Pő+#"[#�U_��[��g� �ET���t-{!��Nr޽�@xy��ww��`�ƍʍ��'�o��V�b�xڼ�������[f����޶m[eP�$$$`Æ�pppDx� �n��ثۇ��B-з�/����vL�lѤY����]_���*�G�������7�
n�>�ȶ�`�_v�#J+]���AV����*��)l�'�����mO-0U3g�q����S;e�H�ۅ:ab��[Ӧ�j�e*�g�u�����r<�@O��;3�����x�x�]��w-�2L8N�:MI�����o�.ZD���]��k�C��OC��M��'�Z�_%
��p*:��01i�}j���q��$^�T����=�u@R�	���E-��kY��v���޽[9:�?�TS1���P�}��,�>�B����ܿ�|uZ�W���ǎV�ăNg��mYY��0��S("�Ԋ٪��z������%mժ5�w�]�~W��k�]#�4���6|�]��16p��`������[$��K�c#��T2J��@I�v�>O���{<�g�n�/�H��."�{���\����s5� �"�.�����
2�᭷ �"�u	R���>]}��]j"@�U����w#Y�z�D�G��i��8��#>�,.%�D~A1؃��H�a���8}�؍F�����6Z��%Eep$�d��eHi��uV��Y���!��a����o�Y��&;g�천�"H4>�g���t�I��*�$�d�� ��J���1�q,�<S}��ot����(4��A�rttt��W#w\�OUjCӌ�m�uD�����+,+F���ѻ���S����>
�>-�}-_̝c�!yю��:.��T�
��j��x�
��'����&r�V���x4k�L!4&:
��|�&_����k�V�|�]wa��G�(�q���x��wT�����x���p��y�_�3g����z��^�	&L��9s�qf,� �6AH���i�^%��{$�#����5_���#r0��(	2L��P��**.ERJ&�X��*Bl�fM��=5�5j42�� %�V���|T��r��V�����Z�"Fe�ܓs��h��Yָp��v��6�#�.[��A�5�7���x�7r)A��@奼�JagS .�Hj��
�󬎙R�x�b��i8�`��@{(��b;9�$6ރE�1%�:΋Q&�fX�5�x!�
�f*�(ъK͈��r�6*��� q�;tζHL�T��q#�������W�PYD�J�iU���Zp�i���f�6E�q�gwn�ۅb��/B��!%bs��DJR��?��PqHf�U�l�TǦw��R:,��[��XP'�$A�j_��y��{j�j+�P�aԻq�iغ�*��j5q�(Z�~6�z�Ze���"�Fo���	�wG��F�b�2�2e��(ր�Aם)&4	$�ի�"��s7�H��^�t����� ��ME��ێ�#���t+��-���nbkY��bkÄᣅ�k�í$�|9��Df����i��Vkj��tx�pWI�u\��������I|p#��yN���*)�uO�[Rf�+@"0���XxE&�0����di��c꤬L�s�������q��sj
�fA�o��=�ܦ ��(G������xe��U�$�܂Y�*
"#A����B7S�T����h���ȹ���R�Z�~�c��AH� tj����|!��_.�llxX �<;1����m5��<�1&=���e|�lG�"Q�~L��*U�˵f����}mhb��;� >$���8�m���#@q��C��[��rS �Ú�7zu��<�nݨ����祦:�:h��"�y �X�X�Td�]9�/�d9�T���KP�77G1�Z��k̞�V�����iu'�����[J��hu��]���D�r\d����,��H�0�ƀh	X/�]6۩۟D#�ۊ� �jX{q��#3�o4R</_��c,�!�^Υ7�� Yx�4���C�5rCA�(]gk��}C굵⮆�u��*���/��4]�^J�jyr�m�K��;���
ь+LN�Ĕ�1U،/��F"[��s\���gmDb[^���S*�i�W[
�s�������3ڴ
$W#G^�ԇ��N��1X�V.ƞ�I}��QF����G���U*5�"�۩v�����p���=|���͙�TD��,^4�"�ɩY��9:ڡM��ծ���A�3r����\߆�~�yy���_���x/7�ұB�I�@q]=T-k��$�����?\����1�a̛�%&OyQͻg^������������ݻ�x�	�7�-�ק#f��"���3ޜ!j׶z�K���~$F;O?����ӄ��С�px���ʜR	RS����[FkhV��R��9"������ ��X��4J�p�	oo�c�}��ܶm;����8��rx�E�^�HT*��ipM�ꄞ%���ԧ�����;1)[wF##������K.���7�"&9�\Bܥ��k#��u���nY�Y����IA�f�|{�*0ผ��i�.mV�AL�|�0bNUy���48�t�w��o���l�L��5#h�1��Qe����_6�������Ho߾Y�2�4/˝f��i�i�
�
�Q<��s�9��QB�*][�!������so�"qdÍ�a���۳�
,9���,[��
��A�^��g�c�~��-�)O���擏?A^���<JĆ�7w�7�9��=�mLM�F��,�Z��A��Ą���]P�BNߗ��ǩ�ީ>��d�*��h��2N��?Kиq�J7ӆde^B���X�ٱ�� S��IL��r�1#��_���ø��{���W7s����<��R�7�1Vvh����B#�ʆ\��+=6�oX�*�u��R3."f򿱖W+*|D�#��h�Q�yz�	7y��UV�QVZ(����`�j]�������Ȕg��MvQ�6�U)��a4|�j�����V�6�������}��L�6YR�����N�~� �ui�%X�`Gu[�^���_c���#A��1?���R4T��,��,�	�v��f�t��܀�Ǐ�d�����7�~Y��/��K/��=��b���ppt���_bݚ���wĠ`ڤ�#[-v�>�+�u�����U��z�s���J�������2x�;�ǽD�B�r"L^��d�Go���*.���Y���,�E��,ą� TTcxMɚ��&�Q�H֊�$�2-q�
K W�ҼyD(:�3���Ғ�1g�/�p�"���"*�v���Bl�0�۽���g륮Y����Vs~���:\QI����캜Եss�~��q~D���H���?�<��O!$4���9+}�P��:�XR[j�˂�:i��Nq{C����˼��J�R)IyΒv�5"��`��n�$ZT7h�����o�X?8=��	��?���z�-����Mj��޽{4	
�������i�	h�OD�BzJ����t'���
��X��+����"�Y78�x�:����P1'������̎��'tv:���)�'����i��\`��"�C�R��ܫ�^`%N�N��4s��	7�3��T/ٝ��Ģ<g̸;7嘷l��Y���.�����+Q[XSA�%�gr�g�������cɒ%��x�r�W�p��Ldeu/u�Li�N�F�ge�D����8	>B!l�3^���M�`����66e��L����=�zR���pE��u�M�(��Y�ZRR��ݏW*cΥ���l���Fj�Z&�>焏T���0�5|:	�&�]1�|�Á�+�0��#(/�߈Ԟ�����jm�,�_@��ͮ2�mZgBX�|��&C��$˪�r�}�D`9t�f��4�����JUYH�p�	ɱq�񙸷L�TU�
��\�MFc�0	�,U+KbM㤔s��u�
gWZ�yM�W2�J���`Mt-�L2�򊣣�MU4Yرڍ�])���vx���b���$�C_Z��g��r��(];E�/(�%�2�q��xx�«�R/'���S��'��N�Қ6m������څ���8WNhպ>��͛#�E[�[��Y��Ĝ0�#t�Y ��K��h�j��o�+��0_c����|GB����5-��<P�A��h������=�E���]��S8�g/��������'����+'��tٹ�'��Αk�Fb���]\�0d��i�_}�U�u�&�����=JT~^.���T\1q�3� �yX�怚4�w�����o�2�����xo���*��i*)�T��`-�é�V-��T�XM����%��c���_|���]�T��u$����}��,v�)lN��7�J�����^z<,���TVO�+d����c��0���p��6*p�BN��Ǳc�Ta��}�nI�O#G���LUpQR���/�(��B���Z��w��{(N�y��L�҄��#�Rk�cNl����$�yRr2�{�9����eZ_/6��I��cɍ�ZBJd��ڌ@��l�p�3<E�pS/9Z���3���L0��a�jH�W��<���P�`�
�nY�aM�5��U毌Ξ�[;G��Fu8q��vK4l���I�G�/V:��%���쐔�������3$m�G�؅ܠF*���!�V��I���ͭߡ]�zl�b>K�+)Q6���t])��b͘���x�M&��h�U|���~\���J�,A'�ԱrPT�N�S5��%$��A�|'�i��I%�ׅ­v�5"�dX���:��ړ323��̨C���)�:���G��,ZrzDTgNN��k�r������|o�^��?5���k�sϷ���@[���Ѯu(��^���+G8떓W��-?"��u���"=�@���;F���kPX����\U�ȅ�߭إ��F��"��ԧ��5�T� .�V���Y�N�w�??�:Eqj6Q�?���&�V@׽!�lP19�s�۬��-#��_��j��z�U�Y�����7v�R�R��L��ET.�l,��(?�̱��go��Á���߫�~�駟��Ύ҉������r}��&�����j�
wm0A~A��s���Or�	�*��m�vGP42ܞ�x����� �r}�g��ևX���TGw�VP���* ��D���XAu9��*�1�\��[W7n�nݺ���t/�$�U�Y�
����O�\r�=1�tÙԼ�����I�D��_�:uR+��.�|��?�\��L��p��~�ݵִ�J�4N�����#�����T\DiZc��F�6A�]����T���{�Y�-]�H���<n]�tQ�
��Âi�B��u�V����� �.*���&L� �'�nE��S�NU'=(�B/�}���\HJ�a$%�618�0L���9h鍞��(-b��Ŋ���O:c�������>Y%٧��Ɔu+�_� �0������cZ�+z�>oo�I��x����k�
� ��n�������Fv��p�āw��E�w�Ġ�Dē�i��w�)Qy>/�C�,|�ll�&�ضm�Z���p!w���i�N�3LIWH�K�6P�F�6�����+*�6*hihC��ZE������+���?�ȑ#��PV	2r�(d^M��}�#�)�$H���Wh!�e�'��������<`���<e�U��o�fa���F�dWX������腶�CP�S��ī8w�r��Еf��{�\J����+�x0�AFb�vϮ���&�] ��6�usjA��ѡm�"���)����l�ZCY�v�3�
j���%���KL���]����,a��E?�l����7q�����99�H���+����#ȠA�����ѵ}ᘊM�γ8]ɸ��"k\��lM�tR��)���s��g:ôd����^��5I�}�]��}�	�W�^�ѭss�s�D����^�8�?��[���n䆗&>��&>%B ��m�XrJ��U��]&ll4Ih����R֌�7���]"�slO�V�?H�b��:k.7�VL/=/����W﹫]H��!X�|��9a���UMe�HNs��_����_o��'�zV���j;+a�9�vm��Ѩc����#뫨B����%���빙K���"�s�V�u�����i��� ���ѻ�a��B������m��-�m|dX�f_}c����������mH��=^��
?_�#��x̹$��]�aC{�i�ojnn����>٫{�%g�%��vi;wǝ}�J��r�D�7�h���#����؞��#F���֫���~>��Ocb��ho��=��io��#N�����=Z-�a{G�����^�r���
C����]>5�L}c�W�>���dCU�b;;�G�K���nuB�RvZ��pC��	�jp���R�P��&z��%G��k����M�v��h�?�b����V�;��H|�pݻ&�����"qe��ٮ.N�T?r�3�ǹ������f����q���P����/5o��D�4q�-\8���U�1b�VH{o3��L�j�͙����CoX��39�XԦ�����l�w��vmB����RDx�&�p���pvTj.�W���h��?���k��M�%�i����3�Th�nE��N�fRq�Fc+u�n弴%���C*Sʹ�47>o��Լ��t��"��.����/n� Qo*@+*UyQ����6U�PEeG���Ș9�}>'R�Z�Le �S�D�Z�;1�7��gÅ�q�tM���j�:J��|L��hm:�6Q5�+����hZs����)8t4���`9��`�NQY��%\'�k�fܘU3^�6/3A`@#5#%�Xno\3�3����I��b	O1U��p�,Ǒ�a����qjr��Dc!�.g�^wvvh�%ƸI���w���e��^D�;ڻ��zl&�
1�R��g�9@�^R�NƉ�i�pm�}��8�?|��,���4�l���+��Z�a�)#�s
|>g�^������G������7|ן��z?-=�OƋ�i���ל+��k3q���A	�36I{G��Q���݈����p��p1��H�g���j+�(Z�2f
Qf	Q>y�)H�6�8H��+,�T�3UKG�����������!�!Kl��K��W��0�ǽ�TVWlJ��M���#9uNM/D��A����ʾ�����7i��o�c�!���@L�F�����S�va/("��X�9��3G�_T����~Q/���p��ȼv#�Du3W�{�ޑA����	bk�_�_OϹC۰��m��>�����:�9���g,7r;y��޸��G$��lu�����`�\�m@\�β�E��pQ�����3�.'��j�9[{W�#�Ï,]�]�����zWR7Oѣ����_X�kpc=]�sR"�Ǧ|$���s	h۩��`�v���/�6�j�Z���l؇�[�T�դ�já�pDeG{Pj}�5`_.�t��8��z�>l�|���ő0�x��=��~ۊ�=�Et�6�J:xќɛ�+�]}۝�>���2t�!��>_���;��v%���&Fp��2�S{WR�<0+99y�h:|<�lX�}{�6�7+��r|b����]{�.�3B�}�D�!�>�M��!�Lz�f`0�[>���g�y{��qٲ�p�l����I�6��V;@$�˜��y���o�}{wG]���O
S{Q
|h�E,���%l����-��g�xl*�l�I��B	�<"��4J����i��: �	��9s�8�f���>�ȹiF�Lo�!����w߭���\0��d&�Rż�j�����r�v�Tտ�&M4�l���Q�8����ȵ�53=3��6¸���3����.������K���N,x�	?˽�s���vi��w�K����:��j�ndn�D!1��#a�0l(A�{�F�ܞ}�v�����/5� �}�ca~���AeR�L���z�!ŵe	S<c�>�6x���n��.6������*G����ݻ�?Y%1�s�6$�J!��x9�GEE�%G ��]��j޼T|蝿��_G`J�aN�\Ȋr�_�����'�u�21�	��](Cf`ތ�D<sW$�-��	�wףp#n���hDDs8:9!'.	�Xi��y����p����EMl���A����̮ݲ4�D�"v.K��Pn[��xIxS%	AD�l3���}���f�ִ����N2��'��	�����C���	i᥼]    IEND�B`�PK   F�X�'  '  /   images/cde853aa-4743-418c-93d3-ccba2bb5bc65.png'�؉PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  &�IDATx��|xT׵�?��z�� 	I� �47�1v(	68�.�7�9��s��9/7��o���;n��8�����P�*�k�5�3��yk�33*����w��u����U���>Ҁ���'����eTT�,l���z����i�������um��	�V��
}[/,VT*n׬V+|}<���
M�]hj�1"����	�iD�ޖ6�h-�=�\�6eB?����#Z��٘_.4�z� 4�<M�h4���Lƞ2:ޠ������`a���K���ha:<ݭ`��4��S�'���U��l��Z����#<��^x��Ό&�Q��I 6zJ�F��	n$-vﻄ�}9x��{��	{
Kj�~���p�NZ�>q��%Z���b�현���>O<F��B[G��;���h��aC˽\�.'�>,$4Ӣ\[d$e]ʿ����+��������!:�AT�����t�J388��%K�����pE{���e/+���e������S'�aD)�7�]t�0�[��.w�X�Է���KO3lAh��O�ۢ��Ѽ�đC�
��X�L�b�|��&��i���c��.?���N�!�Yy���=�{X����u޷Ѳ/o��{�in�Y�n�me����m<7zf�um%X/�Um�3t`Aƽ{��[3�Ͱ��Z���`�6����w�`��LG�����E�F���׊�5�{�������~b��iAyy�x���s6a`�Fd!A�ĝ�@xR<�����8��k� 	�fSA�ރ��kkdL��55u@Mc]�+_G�ƴ��m�,I�T�#���T�o�w�b�V�c��U�o�0��ci�}ro��'��?��R�JׯrCG�A�W �q���Ѹ��i=�����|B��UU��������OO��x�嵰���|�0`�~��d:~����J��A�겏�,?�r%>��(���m�nn.��-��M�����N�߾�*(��$7���KB������(���n��f����U�G�)��94���}FLOJBuu�\���ѳ��F���	_�:z&��֮�RO���У'
���1kv
���c���#����z�4s��ܱc�9����<�b���{!�����,�Դtb��ӡ���'ڌ3��[�a|-Y��MCpP0��dY�V�����(**�G��w8w�E�%K�	O.6��5o�0c�?����
���b��igC ����b�Vqe������ښȊt��Qz~~>1�˗/G||����;s�Z[[�v�Z���)6K����e��'P�'eТ��ׯ_Gzz::��fM�9B��1=1��SH�������^B}c��WSS����ކ�!��4#���CU��h�_/5��������"��ъ/�SCEq8@��� .&��p����Zt>g�UV��	Q�Fy �n����}��@ ��S)�� ύ�ft�����#��2�����F�k,{x�2�5���A8��ϲ�hv�	��nf��7)B�(#8,b2w59�&B�wm?�j#jki�#���$f���0�c��(rk=49otvv�$m6���C�����~>��ҡ��E�5-n�Ї���� �܋S�c�S+�C��@b��� Y����4jn��埭f���	�ۼ6���z/[<ߛ'�v�J(�}���-���E�!���-�/%oЏ7�9��!��ȟ�Ͽ��H����?�!9�Q�ac_#�hd�b��� Ν��ꕙ~�=m�ԳX�IkGT��.�	��MKh���>�n�g��b���Ž�g�esP�`E�{��]�a��5B��<�8jΡ�fΞ=��������⅟�/��V�Ĳ�(���w���|̝3U׫�酻��QX��)����Y�}�b��i��XODGx� Y�ɬCj���u��H���}�o��o,��K Ƅ �`D�ya�]>hhQsCK�_�⃫�f+�
�j��LS�N�@�?04 �CΜ9-AgQf����u���(����s��Hl�7o�%�(--��1������@�J�/AkZ�)�8
��I���.��L���d��U4��`�IyMTԟ��]����sb�����A�_"����o闃�8a	T�PNC�5t͕����t\.k���z>.��y�s�Sŵ�Ƿ�{�ɝ�D�����Ǧ�[ŵ�ܬX����*��G�!1~
��.̜9�Hf���o��O�1C��ǊPXZ��j&R�r�}�.���4Q�$[n:�L��X�M��ݔ�r���H��j@wO�]�r�5��6�����X*k����Jy�AbM��.�6��>�QS�E�@����o���ny�^� � �7�H��F!��V��:�2fK�z�L�$��js
d���x�٧����0>���I(~�U<�%^{�+
���'6��9�j��I����%q����P*kZ�����X��w����C����ڋ�~�-}�����/��K�j)��c�"m�w��=����߿�Gbr+XOXӾή����H�p%�f���[��L�b�c"�-]��R�Ͷ�bE���bǩk�ĉ���[k�����f⅋��w�E�M��W�R�r��t�Y CC&����S��z��^A$V��޽Yҏ���n��=H0�.h��fpt�T���%����� �`'�����ƹB���i+���C>�0i�Q�}�y>Y�����(��C�:
�ވ���[(nE�qǖ'��S�4��@��wv�Ԭ&جF�?{{5S�[�sӹ�/��������	�1e�@��)C��7�k�����.�m�%�;:�U�^��R�W3�1P �;g6f$MGn�%�ڽHII&���ke�����cڴi�Ý�M��=��3䍈)Q�yy'<#�X@]��}���йhp��A��ة"$ψ�#-�g_|�K�ʳ�tM�+��M���b�CF܍��Tf�����E����B�!UWi1���;V{��:��R9�X��J�M��B��d�pZ�C��N��1Է�rýC#�2sz]����9� l�;��h���N�bˆ����������lģ�~�m� ť�Ĭ{���k��%��@жQQQ�q�e�&�fӆ�X�z��:"������ｅ#����/OI&<��+=O}���K \�(O?�����I�B�o��@��@�G��782�@;GU.n��6ː0SE�n�'���y��Z��<¨�s
I$i�����>�,�M��d�|�����b��0okx�hn�v%MHHP�[
APp(����5�ITA����U�Ȫ|s0Yrep�����ic���۪�?������2Y4��o-�!���,�*j�ʠ�d�[HH ڴ� �'�ΟD�%�� �\��˿�wDDƐK$a�5��e�����b�JA2�l�A;SY^�P�|��\����߀b1*z~��Tb]*� �eq�SewK*�r=�`4[a m��V�������v���]Ӽ��kHJJ�+0TC��on������]5����I�s���)G�3�d�9�,�3���q��y��S68d%�r|i�>w�KýK����=��%4ޤ<TG��&�#V�պ���h444`�\���'��<%Oc��
��c Y�J�nR�K�.��\�ncA��ֳ0���d�����i6��!(\ppax�c���&6�3`8/Y�z�Z�������F�v�W�8�c3��b{�da���
���%8�sE�Z�}�*���
�z�nJ(})�4-8� ��Ôq�	J�^�V䴐��6��W�"ƙqhX$f.��(v���3�O����
��H��2�q�d-\�N�P�݅�"
[[��9D�?A�lvAi$����8]�(���	�oh��n��M�Z).�bǯ�+�)������GPP�h���7���8}��\�׷��������oi�=������Fs�D{k�����OBwAeu���A�4�~h=�O���:�7w��X�|>��E�F�����?�qR������p,� YF~�?7K����_�����>����s����w'.���Ծ4��ux��A���|��{b�bAؿ�,*{ wQ\��U��X���aгx�i��zK�(�Ήk�W5cO�b׍8wp��YX_��A���&�"�oR&��P3��ʕb��х�%����!�T��WA5���W��~�J��>��>�y������3�H?.0n��#���� 	LC�~g�y��!���"<M	���}��K|���YgW?N�u��z�$�!!���{`�J�I��T�j���LAY.
��xC	���#��/1GQg�X5�f3*��6��>h��zΦ����N���Ή�+���Lh�����-䭷��)5�,����������$wlhhōF1�s���
7k;�!��0m
��$��F�Gp�|||�:Z^^.4���Ӣa��E�Em?(O�EMn��.9�ze��{��'�g�b	An��c�F\���5J��8"�@�U� �\�3v���R��=v��4>",v��uY���C+2iɓ90��e�������5,.�q���3��"���Px�03~�Ĝ��F�x����=;�5?�LY�g8隔�	^���瀌�=)�N�-��sJ�_�h!���/�Ё�ؾ��-�G�ܙhl�CuM�,JCowN�.�$�qS}�b~�ɮ�V�9�Jb�Z��b�$��3�/�������pP��|� o_>�3\"�4;Q�>$�d��X@l�BSc-����ҷ�)x� ui��K�G��K�R�T�d*8�k6o������D~)
Kj���� -.���q��?JKq�r���-O��u��qqY�fDᅟ>Eq�{���K/����,���8&|��A��B�ł2c.�Yne��v��P�8w�,����o���q�c�����T�[��]�9�;�;	�ċ.��Q�Wä́�J���W�o%{�0P }���`Q�jY%<�*Q�X���=���� ��A֢ę�������/�� ��=��p�5���4i�ܮ�7�����[�p�,��W_%�Svv�q���C�f�v� �t��N-�[�x�u�i�#�w��蘷�X���2�L.0	�Ӎ�H�? f�=�������J�.����a\��(nG���+���� �Ƨ���Im�����:sN�1�:s�"�!��HI�����1h������q�N�Թ)����M߉��H\���-9�ėdb��� &b�Z�
:r�=&0�K�1�M���>2zn�ǎy�kߕ3�Ltaw##.�<��3xl�ZIƸ�544$n�vm�d���!�w�А�ո��y��!�qMJ��� ��ޅҫ�DS�����1�hi�Lln�}�~T�����߈���VQ/1$<���b��Z�R�t-v78s's���x�Br{g�C�k���G�H&�B&� ���NcO'ȍ��a�SP����8�dffJ^�?0H�0
,�ñ�HH�G�|\���ET�<�m�w������L�HY���^�cŊ��{�E���K/�q;Y�s���ٗ�������n� 3nC*�{P~�A�]�#�X�
���Q$����cI)�8a��j��RM���wp�"�!�z����]����r���kp^��f����%�����RF�Ml%��#9y&YN?ZZZ����
�,Ė�N'��x0q]���l9ƶ�Z+������Ϙ�˗������,^8Q�S���{&�V���R�e���ק�8�Z_%.r�'����R�A]�i.�A)�8,DkO�6�8�HO���m������">���Y|{�$�!/$���	���XX�mڄ��p�*�^>-4H���Z�W6�kye;|�#���VW�Efx���Cs�$!u">6Lvj�m�^���-���&dȒ,0^ ��S�̳[���qY%\�t)������,z㾅!���"(��rqQ����/��a�T{��(�Z����r�?T����2ZNq�>�[sh>oV�{���-��[���u)[1�S7��5l��������W˒G��C�CH��;�lQR�WY9s?��1lڸ����;X�r%!��عo��_2&-��\�����������g��p�}8G�ȍ���O��6�U�6�?��0c�=���s�u�Q���W�Y��h����k��$���X�9���V��e�G�n�7D �3$�u]��|�wE�1b"�I��cB�@<hMJJR���*��T�E���^���m��� �'�G�Ɍ��V���l�l��߲e�D�u7����S֥y]{b��ƍj�iq�~?��I��_|IJ9&%�V�����(��Q��+���(�ځS���:'o��D��	B���D��Rb�U����h�7VE(�X�y���8�4V>�=1��^��p���C���k��[ٕ���}��C��|`�<�bf(׿��:)�Tc�ԩ����%A��/n�?1����e�y*�;F(Q\D��s��P���;ضm�Tx9���{�xc^n^>��N�ĵ]=��k2���KIX�|F�.�0PJ!j%��iK�5��ɝ5�&B^�8�XY�陓f&F'y���[���(�1D��S��JA�hjv�-,:�J
�##F<�C�B���OC�_���]Ɯ9s$�O| �h40-&�^z�=f�d���.�V�ܶm[��E �S��s�l³Oo�߿ډ+W�	�
���B��T,��tQ����=v��~���6��ټ��L^k�n�pը�t��\FK��!�b�k׮A��w���sx������x����ąbF=X7twŠ��S4���|Ll���PPP P���H�hf�#�o�v�K�{�hb�6n�(��1O�:%ۂ6oތO>�/^Į=p�RYE���QqwS��G'>\IE?c�k��ǕA�����¢#D��v��&Bg(�;*5��$���&h����&ɜ7�>���j"ƾAsÕ��p��!�����({�fr)�?���Ʋ�b�Ú���J((���2��x|�ܕ����	����@j�0f!�x|�T
X���X��>J:c�]%�ra}NC��D�_�P{�y���fK���J��t�111�ù�D�z��j�Ze�O�cjT����s>�ck[8�J	Ǌ��h�h�)�H&a�	4�,��p_�uܼyS��k�����?�1wӃ}n����p��9����K�a8+ ���&�/�t�����;`� ����/>�^���hқQߤ��xx��wv�fn�\��1I���Q�R�ıYm��c�pcE��kW6�o�&@(����ш��?��(3w��ۈ�n�}�"0�ż
���?�C|BupCY��Qy������K�����Z=	G���:e��^��uyFY��1�����TRBy��
�̓�"���=��Y)F�����k��h�@��Ga�A�c�ю�.E���QRV+��M���x9^�X�r���p�r-!�v<�&����5�����I��N����h��Ƈx��
�O�$�<�+��^{���x��XY[�y���ݱbq4����
q�>X:?� ��,����.]Eiy�n���42
rD \��+%i�����<`1�R|���Nӏ_�x+.�;ػ��ɿ��$�.����݅߿�^��s����cG)L]��g�pa�HP�z����M��c��� �m�ŧ���c�����'ObժUξa�~�=��D�ux]�4܋�2�b��!����",؋r��F��|��Dc� b��,>�σ�͂�H?�X_whMFG��H^���h�+��ᮓk"�}�p�q�ǌ��1�*��}��g��Վݱy�6Vf�{��exhe&4�����a�e��3Y�[�U8s>�*;e�����hn�Ǝ]gP\xQv�\�V�w�y�\�;����Z�AB���p�y077WٰlG�����l/�8���������%u2v�I	X�j9�otK���W������u��<�X07��x����E�� ;� op�1S��u�F=ŋ��N���v|�" q��Xɉ0����q�7gf0	��\����SBQ^�%c(p<'�rT=n/������e�0����O|�mْ��7޼��|��h����?�I�v��R~��*���"e�Vd������F(��j���D���C9��o�8��{"�rrrD ,.rrܺz�*v�9�����7�\(9,-����.I�JJK����!�h�0�����@;Yi[�e7�p�h'a��u��j���Bp[Y:�-7�<z�z`3�p�J�@�~r��a���O�yݽ��lŹ�~�~3:��0@遼�g�V{�tn�R�xa�U�d+nTT4<t�۾�f������"�,5��a������o���`��T�~��5t͚5t~ ���RV�Y�f��SS�L��l�1�w2��U���N)drѲ���`�I�:�7�".�[cs'R�b��N�S3������ȩC().����k)���C/Z��x����&ÅN���ǿDĔp���_}���T�$@R���䋅�\��5�>wݬo��M������5_�E���ܭ�w�8,
�h̷�ٳPUY%[j��f���MG��e�t8]u�����F�f?�OA9�Q+��)֠���'{g�!8��!��M��!+�l1S�ɔ;h2*yÈ᫯�ܴ�+a��p)����Ņ眻y���������J�M�Gn�[��nNMH)1>��&"�ew��P�#�Q���D3��L�?0��(z&�0;?�!� <��
I���(B���M-�&M�hh�Ĭ�L��š����^^�a圛���gNIki�����'��#����XݻBG1�wG4��W�U鷼�梼�6lւ�� ��y0U�>gڮ�@���^9/R-��O�������<M��4���n��d�]�*���y����F��'I��G�j�o?r*����K�#Z���k�볏�s���M����N��oŒ6�3�x���Y1��OX�Ɏ���	���Y޻������*<;�(�~b����w].�Z�����\b��(��z�ǟ��ٟ�|?����ɰ�#��x�f�׮|rWɕ��Y��G�i�3o7�mCցKa\�[�&������E�76|�u4̕��c��Μ�l�墚;�.�UWU��֔Y1����=�r��m��1�{�] W5�z�<�s�+啶��Wڌ�W�r
E��-3#��ֶ�m�3�[��(�1Ԍ�Ľ���m2�,GO	m���{[���2R�-���6/m��[8�%�T�HH�(��&Xf_����)�o�����(�w��*���V�{�3��ڴ9��G�~|mk׶to����-#���ⵇi$ =�6���	x��0��2,�'%�K��YSmY��o�Hퟥ�#�F�m�')����7ζ��Eτ�aBcE�{y<��7/-'ϕm��;4��Et����ϰ�����Ϟ=3�\�o-L���n���`�����8q���W�s*��KM���ג`�y��u,����D��~��1�F�~k��[8���l���f8.�NN�w��m��0�����Wh��k�g̍�w�y��+��5��N�ҏ,(�h�����֜n��c����DS�;�mvZ~a��V��c�үRh���{F��l%L8�`��JN�;���/�/9PF���3���=�b�v��:��Z���S!'ϔ���·٬Ԧ���?M�8h��:�$�J��h_����>%��I�9h#i-��_�cp��Wc�-����9歚�^�� �q4'��j    IEND�B`�PK   F�X�[�"\  o     jsons/user_defined.jsonݖ]o�8��
�5I�m�w,t�h���Eլ��q�6$L>vTU��sB(TJ�ݫ�8���9缯N�ΩS�6{m'6t�ο6��4��C������s����Õ^VkG���2.߬.�m68���st>8��(",6��Oi�������:�@O#���Љ�CCQȕR�����2Rb5C�e��&67Y�*�w�7��gΩ�2�n��e4\k�2�|C����*y�u�8�&QꜾ:I����j�_��v�8	�a��ݏ�w�·W��#*��W	$�pVd1��YV�<���0�%G�R<d��W?���<��vN���SY��V��7�m��M��Dv6��N����'M}��'}��ѧM}V�c�W��������캓ÚZq��k=���M;9��!5w_x����wbDS�:��/e4w�ˆ<?V��U����<��Eoy��y����'�>g��ٳ��mw�5�zw�j�P�F{�Ė�M8���o&���>bw�nB3���DoB�T�-��6)��2��ܒ�x��G�T���e�(�4��CM<���T�Pߏڈ�4��C�:B��`K'�5�c��nNKC�9�c8�5�����v(����g��`(KW6+⍻�X¼��Nm󖫤r�zQVOD�������zN_'�t��Pٻy����n�2��\s�Ʀ�xN'e�MQf6��ݚ�i����a���&Mj�hB�8��e�Q�ae\���5&�$x`��� 'MlR��3��~�)��ڐ.����h�l�7����^���m���4|[�O�� �f�c3��i�7��6���5��[�
d��R�Y��O��if��<t��̃�U�����B`��Mc�I,$js��n�(�aBb��"{��|��z��GkyȼN�#lO�岵>�eo�}���py�/X��f��Т֧���@e:�<�5 ��7�~v~�m�Z�*b�C�!2$��8�:��;n�5 t���c��}�-u��8 �<�w�-�t`Ly6C�𙶘g�{�	�AyLrvH��X�>SrH��������[&�y����c>����h1�[}�1��>�s��]�tm���3��	]�)��(4���ӀD؏$5�n�o PK
   F�X�pǿ�  �C                   cirkitFile.jsonPK
   F�X����V5 GH /             #  images/553717b1-fb1f-43bb-91a8-4009c3c39665.pngPK
   F�Xࢳh� � /             �= images/554ca8bb-9ffd-49bd-8b27-eeb836a64b12.pngPK
   F�X ��ɲ,  �,  /             {� images/c14208cd-713a-4fdc-8661-253b2f19f73c.pngPK
   F�X�'  '  /             z images/cde853aa-4743-418c-93d3-ccba2bb5bc65.pngPK
   F�X�[�"\  o               �D jsons/user_defined.jsonPK      �  sI   